        +          +  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m                                                  "       m  "       m  "       m  "       m  "       m  "       +                                                                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       w  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       m  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�                                                  "       e�  "       e�  "       e�  "       e�  "       e�  "       �                                                                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       �  "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       o  "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       �  "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       e�  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �                                                 "       �p  "       �p  "       �p  "       �p  "       �p  "       �p                                                                                                                          "       �p  "       �p  "       �p  "       �p  "       �p  "       �p              "       �p  "       �p  "       �p                                                                          "       �p  "       �p  "       �p  "       �p  "       �p  "       �p              "       �p  "       �p  "       �p                                                                          "       �p  "       �p  "       �p  "       �p  "       �p  "       �p              "       �p  "       �p                                                                                      "       �p  "       �p  "       �p  "       �p  "       �p  "       �p              "       �p  "       �p  "       �p                                                                          "       �p  "       �p  "       �p  "       �p  "       �p  "       �p              "       �p  "       �p  "       �p                                                                          "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       ~  "       �p  "       �p  "       �p                                                                          "       �p  "       �p  "       �p  "       �p  "       �p  "       �p              "       �p  "       �p                                                                                      "       �p  "       �p  "       �p  "       �p  "       �p  "       �p              "       �p  "       �p                                                                                      "       �p  "       �p  "       �p  "       �p  "       �p  "       �p              "       �p  "       �p  "       �p                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       �p  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`                                                  "       M`  "       M`  "       M`  "       M`  "       M`  "       v                                                                                                                          "       �o  "       �o  "       i`  "       i`  "       �o  "       �o                          "       �o                                                                                      "       l`  "       l`  "       i`  "       i`  "       i`  "       i`              "       o`  "       o`  "       o`                                                                          "       l`  "       l`  "       i`  "       i`  "       i`  "       i`              "       o`  "       o`  "       o`                                                                          "       m`  "       m`  "       j`  "       j`  "       j`  "       j`              "       p`  "       p`  "       p`                                                                          "       m`  "       m`  "       j`  "       j`  "       j`  "       j`              "       p`  "       p`  "       p`                                                                          "       m`  "       m`  "       j`  "       j`  "       j`  "       j`              "       p`  "       p`  "       p`                                                                          "       n`  "       n`  "       k`  "       k`  "       k`  "       k`              "       q`  "       q`                                                                                      "       n`  "       n`  "       k`  "       k`  "       k`  "       k`              "       q`  "       q`                                                                                      "       n`  "       n`  "       k`  "       k`  "       k`  "       k`  "       ?  "       r`  "       q`                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       M`  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,                                                              "       �,  "       �,  "       �,  "       �,  "       �,  "       �,                                                                                                                          "       -  "       -  "       �,  "       �,  "       �,  "       �,              "       -  "       -  "       -                                                                          "       -  "       -  "       �,  "       �,  "       �,  "       �,              "       -  "       -  "       -                                                                          "       -  "       -  "       �,  "       �,  "       �,  "       �,              "       -  "       -  "       -                                                                          "       -  "       -  "       �,  "       �,  "       �,  "       �,              "       -  "       -  "       -                                                                          "       -  "       -  "       �,  "       �,  "       �,  "       �,              "       -  "       -  "       -                                                                          "       -  "       -  "       �,  "       �,  "       �,  "       �,              "       -  "       -  "       -                                                                          "       -  "       -  "        -  "        -  "        -  "        -              "       -  "       -  "       -                                                                          "       -  "       -  "        -  "        -  "        -  "        -              "       -  "       -  "       -                                                                          "       -  "       -  "        -  "        -  "        -  "        -              "       -  "       -  "       -                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       �,  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��                                                  "       ��  "       ��  "       ��  "       ��  "       ��                                                                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                  "       �  "       �  "       �  "       �  "       �                                                                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                              "       �  "       �  "       �  "       �  "       �  "       �                                                                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �          |1          |1  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��                                                  "       ��  "       ��  "       ��  "       ��  "       ��  "       |1                                                                                                                          "       ۳  "       ۳  "       س  "       س  "       س  "       س              "       ޳  "       ޳  "       ޳                                                                          "       ۳  "       ۳  "       س  "       س  "       س  "       س              "       ޳  "       ޳  "       ޳                                                                          "       ۳  "       ۳  "       س  "       س  "       س  "       س  "       m2  "       ޳  "       ޳  "       ޳                                                                          "       ܳ  "       ܳ  "       ٳ  "       ٳ  "       ٳ  "       ٳ              "       ߳  "       ߳                                                                                      "       ܳ  "       ܳ  "       ٳ  "       ٳ  "       ٳ  "       ٳ              "       ߳  "       ߳                                                                                      "       ܳ  "       ܳ  "       ٳ  "       ٳ  "       ٳ  "       ٳ              "       ߳  "       ߳                                                                                      "       ݳ  "       ݳ  "       ڳ  "       ڳ  "       ڳ  "       ڳ                          "       �                                                                                      "       ݳ  "       ݳ  "       ڳ  "       ڳ  "       ڳ  "       ڳ              "       �  "       �                                                                                      "       ݳ  "       ݳ  "       ڳ  "       ڳ  "       ڳ  "       ڳ              "       �  "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S                                                 "       /S "       /S "       /S "       /S "       /S "       "4                                                                                                                          "       NS "       NS "       KS "       KS "       KS "       KS                         "       QS                                                                                     "       NS "       NS "       KS "       KS "       KS "       KS                         "       QS                                                                                     "       NS "       NS "       KS "       KS "       KS "       KS                         "       QS                                                                                     "       OS "       OS "       LS "       LS "       LS "       LS             "       RS "       RS "       RS                                                                         "       OS "       OS "       LS "       LS "       LS "       LS             "       RS "       RS "       RS                                                                         "       OS "       OS "       LS "       LS "       LS "       LS             "       RS "       RS "       RS                                                                         "       PS "       PS "       MS "       MS "       MS "       MS             "       SS "       SS "       SS                                                                         "       PS "       PS "       MS "       MS "       MS "       MS             "       SS "       SS "       SS                                                                         "       PS "       PS "       MS "       MS "       MS "       MS             "       e5  "       SS "       e5                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S "       /S                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:                                                  "       `:  "       `:  "       `:  "       `:  "       `:                                                                                                                                      "       �:  "       �:  "       ~:  "       ~:  "       ~:  "       ~:              "       �:  "       �:                                                                                                              "       ~:  "       ~:                                                                                                                                                  "       �:  "       �:  "       ~:  "       ~:  "       ~:  "       ~:              "       �:  "       �:  "       �:                                                                          "       �:  "       �:  "       :  "       :  "       :  "       :              "       �:  "       �:                                                                                      "       �:  "       �:  "       :  "       :  "       :  "       :              "       �:  "       �:                                                                                      "       �:  "       �:  "       :  "       :  "       :  "       :              "       �:  "       �:  "       �:                                                                          "       �:  "       �:  "       �:  "       �:  "       �:  "       �:              "       �:  "       �:  "       �:                                                                          "       �:  "       �:  "       �:  "       �:  "       �:  "       �:              "       �:  "       �:  "       �:                                                                          "       �:  "       �:  "       �:  "       �:  "       �:  "       �:              "       �:  "       �:  "       �:                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       `:  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       |                                                  "       o  "       o  "       o  "       o  "       o  "       o                                                                                                                          "       s  "       s  "       q  "       q  "       q  "       q              "       v  "       v                                                                                      "       s  "       s  "       q  "       q  "       q  "       q              "       v  "       v  "       v                                                                          "       s  "       s  "       q  "       q  "       q  "       q              "       v  "       v  "       v                                                                          "       t  "       t  "       q  "       q  "       t  "       t              "       w  "       w  "       w                                                                          "       t  "       t  "       q  "       q  "       q  "       q              "       w  "       w  "       w                                                                          "       t  "       t  "       q  "       q  "       q  "       q              "       w  "       w  "       w                                                                          "       u  "       u  "       r  "       r  "       r  "       r              "       x  "       x                                                                                      "       u  "       u  "       r  "       r  "       r  "       r              "       x  "       x                                                                                      "       u  "       u  "       r  "       r  "       r  "       r              "       x  "       x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��                                                  "       ��  "       ��  "       ��  "       ��  "       ��  "       �5                                                                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I                                                 "       I "       I "       I "       I "       I "       �                                                                                                                         "       i "       i "       f "       f "       f "       f             "       l "       l "       l                                                                         "       i "       i "       f "       f "       f "       f             "       l "       l "       l                                                                         "       i "       i "       f "       f "       f "       f             "       l "       l "       l                                                                         "       j "       j "       g "       g "       g "       g             "       m "       m                                                                                     "       j "       j "       g "       g "       g "       g             "       m "       m "       m                                                                         "       j "       j "       g "       g "       g "       g             "       m "       m "       m                                                                         "       k "       k "       h "       h "       h "       h             "       n "       n "       n                                                                         "       k "       k "       h "       h "       h "       h             "       n "       n                                                                                     "       k "       k "       h "       h "       h "       h             "       n "       n "       n                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I "       I         �          �  "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "                                                         "         "         "         "         "         "       �                                                                                                                          "       #  "       #  "          "          "          "                      "       &  "       &  "       &                                                                          "       #  "       #  "          "          "          "                      "       &  "       &  "       &                                                                          "       #  "       #  "          "          "          "                      "       &  "       &                                                                                      "       $  "       $  "       !  "       !  "       !  "       !              "       '  "       '  "       '                                                                          "       $  "       $  "       !  "       !  "       !  "       !              "       '  "       '  "       '                                                                          "       $  "       $  "       !  "       !  "       !  "       !              "       '  "       '                                                                                      "       %  "       %  "       "  "       "  "       "  "       "                          "       (                                                                                      "       %  "       %  "       "  "       "  "       "  "       "              "       (  "       (  "       (                                                                          "       %  "       %  "       "  "       "  "       "  "       "              "       (  "       (  "       (                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "         "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��                                                  "       ��  "       ��  "       ��  "       ��  "       ��  "       �5                                                                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��                                                                                                              "       ��  "       ��                                                                                                                                                  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       Zb                                                 "       � "       � "       � "       � "       � "       �                                                                                                                         "       � "       � "       � "       � "       � "       �             "       � "       � "       �                                                                         "       � "       � "       � "       � "       � "       �             "       � "       �                                                                                     "       � "       � "       � "       � "       � "       �             "       � "       �                                                                                     "       � "       � "       � "       � "       � "       �             "       � "       � "       �                                                                         "       � "       � "       � "       � "       � "       �             "       � "       � "       �                                                                         "       � "       � "       � "       � "       � "       �             "       � "       � "       �                                                                         "       � "       � "       � "       � "       � "       �             "       � "       � "       �                                                                         "       � "       � "       � "       � "       � "       �             "       � "       � "       �                                                                         "       � "       � "       � "       � "       � "       �             "       � "       � "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A                                                  "       A  "       A  "       A  "       A  "       A                                                                                                                                      "       `  "       `  "       ]  "       ]  "       ]  "       ]              "       c  "       c                                                                                      "       `  "       `  "       ]  "       ]  "       ]  "       ]              "       c  "       c  "       c                                                                          "       `  "       `  "       ]  "       ]  "       ]  "       ]              "       c  "       c  "       c                                                                          "       a  "       a  "       ^  "       ^  "       ^  "       ^              "       d  "       d  "       d                                                                          "       a  "       a  "       ^  "       ^  "       ^  "       ^              "       d  "       d  "       d                                                                          "       a  "       a  "       ^  "       ^  "       ^  "       ^              "       d  "       d                                                                                      "       b  "       b  "       _  "       _  "       _  "       _              "       e  "       e  "       e                                                                          "       b  "       b  "       _  "       _  "       _  "       _              "       e  "       e                                                                                      "       b  "       b  "       _  "       _  "       _  "       _              "       e  "       e  "       e                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A                                                  "       �A  "       �A  "       �A  "       �A  "       �A  "       �                                                                                                                          "       B  "       B  "       B  "       B  "       B  "       B              "       B  "       B  "       B                                                                          "       B  "       B  "       B  "       B  "       B  "       B              "       B  "       B  "       B                                                                          "       B  "       B  "       B  "       B  "       B  "       B              "       B  "       B  "       B                                                                          "       B  "       B  "       B  "       B  "       B  "       B              "       B  "       B  "       B                                                                          "       B  "       B  "       B  "       B  "       B  "       B              "       B  "       B  "       B                                                                          "       B  "       B  "       B  "       B  "       B  "       B              "       B  "       B  "       B                                                                          "       B  "       B  "       B  "       B  "       B  "       B              "       B  "       B  "       B                                                                          "       B  "       B  "       B  "       B  "       B  "       B              "       B  "       B  "       B                                                                          "       B  "       B  "       B  "       B  "       B  "       B              "       B  "       B  "       B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �A  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7                                                              "       �7  "       �7  "       �7  "       �7  "       �7  "       �7                                                                                                                          "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7  "       �7                                                                          "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7  "       �7                                                                          "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7  "       �7                                                                          "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7                                                                                      "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7                                                                                      "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7  "       �7                                                                          "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7                                                                                      "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7                                                                                      "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c                                                             "       c "       c "       c "       c "       c "       c                                                                                                                         "       c "       c "       c "       c "       c "       c                         "       c                                                                                     "       c "       c "       c "       c "       c "       c                         "       c                                                                                     "       c "       c "       c "       c "       c "       c                         "       c                                                                                     "       c "       c "       c "       c "       c "       c             "       c "       c "       c                                                                         "       c "       c "       c "       c "       c "       c             "       c "       c "       c                                                                         "       c "       c "       c "       c "       c "       c                         "       c                                                                                     "       c "       c "       c "       c "       c "       c             "       c "       c "       c                                                                         "       c "       c "       c "       c "       c "       c             "       c "       c                                                                                     "       c "       c "       c "       c "       c "       c             "       c "       c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c "       c                   "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "                                                        "       �  "       �  "       �  "       �  "       �  "       �                                                                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                                              "       �  "       �                                                                                                                                                  "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6                                                  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6                                                                                                                          "       �6  "       �6  "       �6  "       �6  "       �6  "       �6              "       �6  "       �6  "       �6                                                                          "       �6  "       �6  "       �6  "       �6  "       �6  "       �6              "       �6  "       �6                                                                                      "       �6  "       �6  "       �6  "       �6  "       �6  "       �6              "       �6  "       �6                                                                                      "       �6  "       �6  "       �6  "       �6  "       �6  "       �6              "       �6  "       �6                                                                                      "       �6  "       �6  "       �6  "       �6  "       �6  "       �6              "       �6  "       �6                                                                                      "       �6  "       �6  "       �6  "       �6  "       �6  "       �6              "       �6  "       �6  "       �6                                                                          "       �6  "       �6  "       �6  "       �6  "       �6  "       �6              "       �6  "       �6  "       �6                                                                          "       �6  "       �6  "       �6  "       �6  "       �6  "       �6              "       �6  "       �6  "       �6                                                                          "       �6  "       �6  "       �6  "       �6  "       �6  "       �6              "       �6  "       �6  "       �6                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       �6  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7                                                              "       :7  "       :7  "       :7  "       :7  "       :7  "       :7                                                                                                                          "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7                                                                                      "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7                                                                                      "       �7  "       �7  "       �7  "       �7  "       �7  "       �7  "       2O  "       �7  "       �7  "       �7                                                                          "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7  "       �7                                                                          "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7  "       �7                                                                          "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7  "       �7                                                                          "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7                                                                                      "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7  "       �7                                                                          "       �7  "       �7  "       �7  "       �7  "       �7  "       �7              "       �7  "       �7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       :7  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#                                                  "       �#  "       �#  "       �#  "       �#  "       �#                                                                                                                                      "       �#  "       �#  "       �#  "       �#  "       �#  "       �#              "       �#  "       �#  "       �#                                                                          "       �#  "       �#  "       �#  "       �#  "       �#  "       �#              "       �#  "       �#  "       �#                                                                          "       �#  "       �#  "       �#  "       �#  "       �#  "       �#              "       �#  "       �#  "       �#                                                                          "       �#  "       �#  "       �#  "       �#  "       �#  "       �#              "       �#  "       �#                                                                                      "       �#  "       �#  "       �#  "       �#  "       �#  "       �#              "       �#  "       �#  "       �#                                                                          "       �#  "       �#  "       �#  "       �#  "       �#  "       �#              "       �#  "       �#  "       �#                                                                          "       �#  "       �#  "       �#  "       �#  "       �#  "       �#              "       �#  "       �#  "       �#                                                                          "       �#  "       �#  "       �#  "       �#  "       �#  "       �#              "       �#  "       �#  "       �#                                                                          "       �#  "       �#  "       �#  "       �#  "       �#  "       �#              "       �#  "       �#  "       �#                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[                                                              "       �[  "       �[  "       �[  "       �[  "       �[  "       �[                                                                                                                          "       �[  "       �[  "       �[  "       �[  "       �[  "       �[              "       �[  "       �[  "       �[                                                                          "       �[  "       �[  "       �[  "       �[  "       �[  "       �[              "       �[  "       �[  "       �[                                                                          "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �m  "       �[  "       �[  "       �[                                                                          "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �g  "       Fg  "       �[  "       Fg                                                                          "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       o  "       �[  "       �[  "       �[                                                                          "       �[  "       �[  "       �[  "       �[  "       �[  "       �[              "       �[  "       �[  "       �[                                                                          "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �e  "       e  "       �[  "       e                                                                          "       �[  "       �[  "       �[  "       �[  "       �[  "       �[                          "       �[                                                                                      "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       d  "       �[  "       �[  "       �[                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[  "       �[                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �%                                                 "       �% "       �% "       �% "       �% "       �%                                                                                                                                     "       �% "       �% "       �% "       �% "       �% "       �%             "       �% "       �% "       �%                                                                         "       �% "       �% "       �% "       �% "       �% "       �%             "       �% "       �%                                                                                     "       �% "       �% "       �% "       �% "       �% "       �%             "       �% "       �%                                                                                     "       �% "       �% "       �% "       �% "       �% "       �%             "       �% "       �% "       �%                                                                         "       �% "       �% "       �% "       �% "       �% "       �%             "       �% "       �% "       �%                                                                         "       �% "       �% "       �% "       �% "       �% "       �%             "       �% "       �% "       �%                                                                         "       �% "       �% "       �% "       �% "       �% "       �%             "       �% "       �% "       �%                                                                         "       �% "       �% "       �% "       �% "       �% "       �%             "       �% "       �%                                                                                     "       �% "       �% "       �% "       �% "       �% "       �%             "       �% "       �%                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �% "       �%         Ѝ          Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ                                                  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ                                                                                                                                      "       ��  "       ��  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       ��  "       ��  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       ��  "       ��  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �                          "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �                          "       ��                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       ��  "       ��  "       ��                                                                          "       �  "       �  "       �  "       �  "       �  "       �                          "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Ѝ  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv                                                              "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv                                                                                                                          "       Gv  "       Gv  "       Ev  "       Ev  "       Ev  "       Ev              "       Jv  "       Jv  "       Jv                                                                          "       Gv  "       Gv  "       Ev  "       Ev  "       Ev  "       Ev              "       Jv  "       Jv  "       Jv                                                                          "       Gv  "       Gv  "       Ev  "       Ev  "       Ev  "       Ev              "       Jv  "       Jv  "       Jv                                                                          "       Hv  "       Hv  "       Ev  "       Ev  "       Ev  "       Ev              "       Kv  "       Kv  "       Kv                                                                          "       Hv  "       Hv  "       Ev  "       Ev  "       Ev  "       Ev              "       Kv  "       Kv  "       Kv                                                                          "       Hv  "       Hv  "       Ev  "       Ev  "       Ev  "       Ev              "       Kv  "       Kv                                                                                      "       Iv  "       Iv  "       Fv  "       Fv  "       Fv  "       Fv              "       Lv  "       Lv  "       Lv                                                                          "       Iv  "       Iv  "       Fv  "       Fv  "       Fv  "       Fv              "       Lv  "       Lv  "       Lv                                                                          "       Iv  "       Iv  "       Fv  "       Fv  "       Fv  "       Fv              "       Mv  "       Lv  "       Lv                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       Cv  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�                                                  "       }�  "       }�  "       }�  "       }�  "       }�                                                                                                                                      "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       j "       j "       ��  "       ��  "       j "       j             "       j "       j "       j                                                                         "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                                                  "       ��  "       ��                                                                                                                                                                          "       ��  "       ��                                                                                                                                                  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��              "       ��  "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       }�  "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E&                                                             "       E& "       E& "       E& "       E& "       E& "       E&                                                                                                                         "       I& "       I& "       G& "       G& "       G& "       G&             "       L& "       L&                                                                                     "       I& "       I& "       G& "       G& "       G& "       G&             "       L& "       L& "       L&                                                                         "       I& "       I& "       G& "       G& "       G& "       G&             "       L& "       L& "       L&                                                                         "       J& "       J& "       G& "       G& "       G& "       G&             "       M& "       M&                                                                                     "       J& "       J& "       G& "       G& "       G& "       G&             "       M& "       M& "       M&                                                                         "       J& "       J& "       G& "       G& "       G& "       G&             "       M& "       M&                                                                                     "       K& "       K& "       H& "       H& "       H& "       H&             "       N& "       N&                                                                                     "       K& "       K& "       H& "       H& "       H& "       H&             "       N& "       N&                                                                                     "       K& "       K& "       H& "       H& "       H& "       H&             "       N& "       N&                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E& "       E&                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��                                                  "       ��  "       ��  "       ��  "       ��  "       ��  "       pt                                                                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       ]y  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       �{  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       �v  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       x  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �  "       |  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                  "       �  "       �  "       �  "       �  "       �  "       �~                                                                                                                          "       =�  "       =�  "       :�  "       :�  "       :�  "       :�              "       @�  "       @�  "       @�                                                                          "       =�  "       =�  "       :�  "       :�  "       :�  "       :�              "       @�  "       @�  "       @�                                                                          "       =�  "       =�  "       :�  "       :�  "       :�  "       :�              "       @�  "       @�  "       @�                                                                          "       >�  "       >�  "       ;�  "       ;�  "       ;�  "       ;�              "       A�  "       A�  "       A�                                                                          "       >�  "       >�  "       ;�  "       ;�  "       ;�  "       ;�              "       A�  "       A�  "       A�                                                                          "       >�  "       >�  "       ;�  "       ;�  "       ;�  "       ;�              "       A�  "       A�  "       A�                                                                          "       ?�  "       ?�  "       <�  "       <�  "       <�  "       <�              "       B�  "       B�  "       B�                                                                          "       ?�  "       ?�  "       <�  "       <�  "       <�  "       <�              "       B�  "       B�  "       B�                                                                          "       ?�  "       ?�  "       <�  "       <�  "       <�  "       <�              "       B�  "       B�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                              "       �  "       �  "       �  "       �  "       �  "       �                                                                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       :�  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       ]�  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       *�  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �  "       $�  "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��                                                              "       ��  "       ��  "       ��  "       ��  "       ��  "       ��                                                                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       �  "       �  "       �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "        �  "        �  "        �                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       4�  "        �  "       4�                                                                                                  "       �  "       �                                                                                                                                                  "       �  "       �  "       �  "       �  "       �  "       �              "       !�  "       !�  "       !�                                                                          "       �  "       �  "       �  "       �  "       �  "       �              "       !�  "       !�                                                                                      "       �  "       �  "       �  "       �  "       �  "       �              "       !�  "       !�  "       !�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+                                                  "       3+  "       3+  "       3+  "       3+  "       3+                                                                                                                                      "       R+  "       R+  "       O+  "       O+  "       O+  "       O+                          "       U+                                                                                      "       R+  "       R+  "       O+  "       O+  "       O+  "       O+              "       U+  "       U+  "       U+                                                                          "       R+  "       R+  "       O+  "       O+  "       O+  "       O+              "       U+  "       U+  "       U+                                                                          "       S+  "       S+  "       P+  "       P+  "       P+  "       P+              "       V+  "       V+  "       V+                                                                          "       S+  "       S+  "       P+  "       P+  "       P+  "       P+              "       V+  "       V+  "       V+                                                                          "       S+  "       S+  "       P+  "       P+  "       P+  "       P+              "       V+  "       V+  "       V+                                                                          "       T+  "       T+  "       Q+  "       Q+  "       Q+  "       Q+              "       W+  "       W+                                                                                      "       T+  "       T+  "       Q+  "       Q+  "       Q+  "       Q+              "       W+  "       W+                                                                                      "       T+  "       T+  "       Q+  "       Q+  "       Q+  "       Q+              "       X+  "       W+  "       W+                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+  "       3+                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�                                                  "       &�  "       &�  "       &�  "       &�  "       &�                                                                                                                                      "       F�  "       F�  "       C�  "       C�  "       C�  "       C�              "       I�  "       I�  "       I�                                                                          "       F�  "       F�  "       C�  "       C�  "       C�  "       C�              "       I�  "       I�  "       I�                                                                          "       ��  "       ��  "       C�  "       C�  "       ��  "       ��              "       ��  "       ��  "       ��                                                                          "       G�  "       G�  "       D�  "       D�  "       D�  "       D�                          "       J�                                                                                      "       G�  "       G�  "       D�  "       D�  "       D�  "       D�                          "       J�                                                                                      "       G�  "       G�  "       D�  "       D�  "       D�  "       D�                          "       J�                                                                                      "       H�  "       H�  "       E�  "       E�  "       E�  "       E�                          "       K�                                                                                      "       H�  "       H�  "       E�  "       E�  "       E�  "       E�                          "       K�                                                                                      "       H�  "       H�  "       E�  "       E�  "       E�  "       E�              "       K�  "       K�  "       K�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       &�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�                                                              "       E�  "       E�  "       E�  "       E�  "       E�  "       E�                                                                                                                          "       I�  "       I�  "       G�  "       G�  "       G�  "       G�              "       L�  "       L�                                                                                      "       I�  "       I�  "       G�  "       G�  "       G�  "       G�              "       L�  "       L�                                                                                      "       I�  "       I�  "       G�  "       G�  "       G�  "       G�              "       L�  "       L�                                                                                      "       J�  "       J�  "       G�  "       G�  "       G�  "       G�              "       M�  "       M�  "       M�                                                                          "       J�  "       J�  "       G�  "       G�  "       G�  "       G�              "       M�  "       M�  "       M�                                                                          "       J�  "       J�  "       G�  "       G�  "       G�  "       G�              "       M�  "       M�  "       M�                                                                          "       K�  "       K�  "       H�  "       H�  "       H�  "       H�              "       N�  "       N�  "       N�                                                                          "       K�  "       K�  "       H�  "       H�  "       H�  "       H�              "       N�  "       N�  "       N�                                                                          "       K�  "       K�  "       H�  "       H�  "       H�  "       H�              "       N�  "       N�  "       N�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�  "       E�          D         D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D                                                 "       D "       D "       D "       D "       D                                                                                                                                     "       !D "       !D "       D "       D "       D "       D             "       $D "       $D "       $D                                                                         "       !D "       !D "       D "       D "       D "       D             "       $D "       $D "       $D                                                                         "       !D "       !D "       D "       D "       D "       D             "       $D "       $D                                                                                     "       "D "       "D "       D "       D "       D "       D             "       %D "       %D                                                                                     "       "D "       "D "       D "       D "       D "       D             "       %D "       %D                                                                                     "       "D "       "D "       D "       D "       D "       D             "       %D "       %D                                                                                     "       #D "       #D "        D "        D "        D "        D             "       &D "       &D "       &D                                                                         "       #D "       #D "        D "        D "        D "        D             "       &D "       &D "       &D                                                                         "       #D "       #D "        D "        D "        D "        D             "       &D "       &D "       &D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D "       D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�                                                  "       R�  "       R�  "       R�  "       R�  "       R�  "       ��                                                                                                                          "       s�  "       s�  "       p�  "       p�  "       p�  "       p�              "       v�  "       v�  "       v�                                                                          "       s�  "       s�  "       p�  "       p�  "       p�  "       p�              "       v�  "       v�  "       v�                                                                          "       s�  "       s�  "       p�  "       p�  "       p�  "       p�              "       v�  "       v�  "       v�                                                                                                  "       q�  "       q�                                                                                                                                                  "       t�  "       t�  "       q�  "       q�  "       q�  "       q�              "       w�  "       w�  "       w�                                                                          "       t�  "       t�  "       q�  "       q�  "       q�  "       q�              "       w�  "       w�  "       w�                                                                          "       u�  "       u�  "       r�  "       r�  "       r�  "       r�              "       x�  "       x�  "       x�                                                                          "       u�  "       u�  "       r�  "       r�  "       r�  "       r�  "       g�  "       x�  "       x�  "       x�                                                                          "       u�  "       u�  "       r�  "       r�  "       r�  "       r�              "       x�  "       x�  "       x�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�                                                              "       N�  "       N�  "       N�  "       N�  "       N�  "       N�                                                                                                                                                  "       ��  "       ��  "       ��  "       ��                                                                                                                                                  "       ��  "       ��  "       ��  "       ��                                                                                                                                                  "       ��  "       ��  "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       N�  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w                                                  "       w  "       w  "       w  "       w  "       w                                                                                                                                      "       .w  "       .w  "       +w  "       +w  "       +w  "       +w              "       1w  "       1w                                                                                      "       .w  "       .w  "       +w  "       +w  "       +w  "       +w              "       1w  "       1w                                                                                      "       .w  "       .w  "       +w  "       +w  "       +w  "       +w              "       1w  "       1w                                                                                      "       /w  "       /w  "       ,w  "       ,w  "       ,w  "       ,w              "       2w  "       2w                                                                                      "       /w  "       /w  "       ,w  "       ,w  "       ,w  "       ,w              "       2w  "       2w                                                                                      "       /w  "       /w  "       ,w  "       ,w  "       ,w  "       ,w              "       2w  "       2w                                                                                      "       0w  "       0w  "       -w  "       -w  "       -w  "       -w              "       3w  "       3w                                                                                      "       0w  "       0w  "       -w  "       -w  "       -w  "       -w              "       3w  "       3w  "       3w                                                                          "       0w  "       0w  "       -w  "       -w  "       -w  "       -w              "       3w  "       3w  "       3w                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       w  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       ��                                                  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx                                                                                                                          "       �x  "       �x  "       �x  "       �x  "       �x  "       �x                          "       �x                                                                                      "       �x  "       �x  "       �x  "       �x  "       �x  "       �x                          "       �x                                                                                      "       �x  "       �x  "       �x  "       �x  "       �x  "       �x              "       �x  "       �x                                                                                      "       �x  "       �x  "       �x  "       �x  "       �x  "       �x                          "       �x                                                                                      "       �x  "       �x  "       �x  "       �x  "       �x  "       �x              "       �x  "       �x                                                                                      "       �x  "       �x  "       �x  "       �x  "       �x  "       �x              "       �x  "       �x  "       �x                                                                          "       �x  "       �x  "       �x  "       �x  "       �x  "       �x              "       �x  "       �x  "       �x                                                                          "       �x  "       �x  "       �x  "       �x  "       �x  "       �x              "       �x  "       �x  "       �x                                                                          "       �x  "       �x  "       �x  "       �x  "       �x  "       �x              "       �x  "       �x                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx  "       xx                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          :�          :�  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X                                                  "       �X  "       �X  "       �X  "       �X  "       �X                                                                                                                                      "       �X  "       �X  "       �X  "       �X  "       �X  "       �X              "       �X  "       �X  "       �X                                                                          "       �X  "       �X  "       �X  "       �X  "       �X  "       �X              "       �X  "       �X                                                                                      "       �X  "       �X  "       �X  "       �X  "       �X  "       �X              "       �X  "       �X  "       �X                                                                          "       �X  "       �X  "       �X  "       �X  "       �X  "       �X              "       �X  "       �X                                                                                      "       �X  "       �X  "       �X  "       �X  "       �X  "       �X              "       �X  "       �X                                                                                      "       �X  "       �X  "       �X  "       �X  "       �X  "       �X              "       �X  "       �X                                                                                      "       �X  "       �X  "       �X  "       �X  "       �X  "       �X              "       �X  "       �X  "       �X                                                                          "       �X  "       �X  "       �X  "       �X  "       �X  "       �X              "       �X  "       �X  "       �X                                                                          "       �X  "       �X  "       �X  "       �X  "       �X  "       �X              "       �X  "       �X  "       �X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X  "       �X                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g                                                  "       �g  "       �g  "       �g  "       �g  "       �g                                                                                                                                                              "       �g  "       �g                                                                                                                                                                          "       �g  "       �g                                                                                                                                                  "       h  "       h  "       �g  "       �g  "       �g  "       �g              "       h  "       h  "       h                                                                          "       h  "       h  "        h  "        h  "        h  "        h              "       h  "       h  "       h                                                                          "       h  "       h  "        h  "        h  "        h  "        h              "       h  "       h  "       h                                                                          "       h  "       h  "        h  "        h  "        h  "        h              "       h  "       h  "       h                                                                          "       h  "       h  "       h  "       h  "       h  "       h              "       h  "       h  "       h                                                                          "       h  "       h  "       h  "       h  "       h  "       h              "       h  "       h  "       h                                                                          "       h  "       h  "       h  "       h  "       h  "       h  "       Ci  "       h  "       h  "       h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       �g  "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       �                                                 "       � "       � "       � "       � "       �                                                                                                                                     "       � "       � "       � "       � "       � "       �             "       � "       �                                                                                     "       � "       � "       � "       � "       � "       �             "       � "       �                                                                                     "       � "       � "       � "       � "       � "       �             "       � "       �                                                                                     "       � "       � "       � "       � "       � "       �             "       � "       � "       �                                                                         "       � "       � "       � "       � "       � "       �             "       � "       � "       �                                                                         "       � "       � "       � "       � "       � "       �             "       � "       � "       �                                                                         "       � "       � "       � "       � "       � "       �             "       � "       � "       �                                                                         "       � "       � "       � "       � "       � "       �             "       � "       �                                                                                     "       � "       � "       � "       � "       � "       �             "       � "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       � "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �~                                                  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I                                                                                                                          "       J  "       J  "       J  "       J  "       J  "       J                          "       J                                                                                      "       J  "       J  "       J  "       J  "       J  "       J                          "       J                                                                                      "       J  "       J  "       J  "       J  "       J  "       J                          "       J                                                                                      "       J  "       J  "       J  "       J  "       J  "       J              "       J  "       J  "       J                                                                          "       J  "       J  "       J  "       J  "       J  "       J              "       J  "       J  "       J                                                                          "       J  "       J  "       J  "       J  "       J  "       J              "       J  "       J                                                                                      "       J  "       J  "       J  "       J  "       J  "       J              "       J  "       J  "       J                                                                          "       J  "       J  "       J  "       J  "       J  "       J              "       J  "       J                                                                                      "       J  "       J  "       J  "       J  "       J  "       J              "       J  "       J  "       J                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I                                                  "       �I  "       �I  "       �I  "       �I  "       �I  "       /J                                                                                                                          "       �I  "       �I  "       �I  "       �I  "       �I  "       �I                          "       �I                                                                                      "       �I  "       �I  "       �I  "       �I  "       �I  "       �I              "       �I  "       �I  "       �I                                                                          "       �I  "       �I  "       �I  "       �I  "       �I  "       �I              "       �I  "       �I  "       �I                                                                          "       �I  "       �I  "       �I  "       �I  "       �I  "       �I              "       �I  "       �I                                                                                      "       �I  "       �I  "       �I  "       �I  "       �I  "       �I              "       �I  "       �I                                                                                      "       �I  "       �I  "       �I  "       �I  "       �I  "       �I              "       �I  "       �I  "       �I                                                                          "       �I  "       �I  "       �I  "       �I  "       �I  "       �I              "       �I  "       �I  "       �I                                                                          "       �I  "       �I  "       �I  "       �I  "       �I  "       �I              "       �I  "       �I  "       �I                                                                          "       �I  "       �I  "       �I  "       �I  "       �I  "       �I              "       �I  "       �I  "       �I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       ]�  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       ^�  "       ^�  "       ^�  "       ^�  "       �D  "       ^�  "       ^�  "       ^�  "       ^�  "       �D  "       �D  "       �D  "       �D  "       �D  "       ^�  "       ^�  "       ^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �#  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       <  "       <  "       <  "       <  "       <  "       <  "       <  "       <  "       <  "       <  "       <  "       <  "       =  "       =  "       =  "       =  "       =  "       =  "       =  "       =  "       =  "       =  "       =  "       =  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       ?  "       ?  "       ?  "       ?  "       ?  "       ?  "       ?  "       ?  "       ?  "       ?  "       ?  "       ?  "       @  "       @  "       @  "       @  "       @  "       @  "       @  "       @  "       @  "       @  "       @  "       @  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       A  "       B  "       B  "       B  "       B  "       B  "       B  "       B  "       B  "       B  "       B  "       B  "       B  "       C  "       C  "       C  "       C  "       C  "       C  "       C  "       C  "       C  "       C  "       C  "       C  "       D  "       D  "       D  "       D  "       D  "       D  "       D  "       D  "       D  "       D  "       D  "       D  "       E  "       E  "       E  "       E  "       E  "       E  "       E  "       E  "       E  "       E  "       E  "       E  "       F  "       F  "       F  "       F  "       F  "       F  "       F  "       F  "       F  "       F  "       F  "       F  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       H  "       H  "       H  "       H  "       H  "       H  "       H  "       H  "       H  "       H  "       H  "       H  "       I  "       I  "       I  "       I  "       I  "       I  "       I  "       I  "       I  "       I  "       I  "       I  "       �   "       �   "       �   "       �   "       �   "       �   "       �                                                   "       �                                                   "       �   "       �   "       �   "       �   "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       9  "       9  "       9  "       9  "       9  "       9  "       9                                                  "       9                                                  "       9  "       9  "       9  "       9  "       9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       9  "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �                                                   "       �                                                   "       �   "       �   "       �   "       �   "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   &       n  &       n  &       n  &       n  &         &         &         &         &       O`  &       O`  &       O`  &       O`  &       N`  &       N`  &       N`  &       N`  &         &         &         &         &         &         &         &         &       +�  &       +�  &       +�  &       +�  &       �+  &       �+  &       �+  &       �+  &       O`  &       O`  &       O`  &       O`  &         &         &         &         &         &         &         &         &         &         &         &         &       4+  &       4+  &       4+  &       4+  &       4+  &       4+  &       4+  &       4+  &       n  &       n  &       n  &       n  &       n  &       n  &       n  &       n  &       n  &       n  &       n  &       n                                                  &       o  &       o  &       o  &       o                                                  &       ��  &       ��  &       ��  &       ��                                                  &         &         &         &         &       zo  &       zo  &       zo  &       zo  &         &         &         &         &       N`  &       N`  &       N`  &       N`  &       N`  &       N`  &       N`  &       N`  &         &         &         &         &       N`  &       N`  &       N`  &       N`  &       �`  &       �`  &       �`  &       �`  &       n  &       n  &       n  &       n  &       4+  &       4+  &       4+  &       4+  &       4+  &       4+  &       4+  &       4+  &       4+  &       4+  &       4+  &       4+  &       n  &       n  &       n  &       n  &       4+  &       4+  &       4+  &       4+  &       o  &       o  &       o  &       o  &         &         &         &         &       O`  &       O`  &       O`  &       O`  &       O`  &       O`  &       O`  &       O`  &       n  &       n  &       n  &       n  &       n  &       n  &       n  &       n                                                  &       N`  &       N`  &       N`  &       N`  &       n  &       n  &       n  &       n  &       O`  &       O`  &       O`  &       O`  &       O`  &       O`  &       O`  &       O`  &       n  &       n  &       n  &       n  &         &         &         &         &       ҍ  &       ҍ  &       ҍ  &       ҍ  &       S  &       S  &       S  &       S  &       �  &       �  &       �  &       �  &       ��  &       ��  &       ��  &       ��  &       �@  &       �@  &       �@  &       �@  &       o  &       o  &       o  &       o  &       o  &       o  &       o  &       o  &       S  &       S  &       S  &       S  &       ��  &       ��  &       ��  &       ��  &       D &       D &       D &       D &       4+  &       4+  &       4+  &       4+  &       n  &       n  &       n  &       n  &       n  &       n  &       n  &       o  &       n  &       n  &       n  &       n  &       �V  &       �V  &       �V  &       �V  &       �  &       �  &       �  &       �  &       �X  &       �X  &       �X  &       �X  &       D- &       D- &       D- &       D- &       D- &       D- &       D- &       D- &       �X  &       �X  &       �X  &       �X  &       KZ  &       KZ  &       KZ  &       KZ                                                                                                  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �X  &       �X  &       �X  &       �X  &       b�  &       b�  &       b�  &       b�  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �                                                  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �X  &       �X  &       �X  &       �X  &       �X  &       �X  &       �X  &       �X  &       �:  &       �:  &       �:  &       �:  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �                                                  &       �  &       �  &       �  &       �  &       �X  &       �X  &       �X  &       �X  &       �:  &       �:  &       �:  &       �:  &       �X  &       �X  &       �X  &       �X  &       �X  &       �X  &       �X  &       �X  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �X  &       �X  &       �X  &       �X  &       �,  &       �,  &       �,  &       �,                                                  &       +Z  &       +Z  &       +Z  &       +Z  &       ;Z  &       ;Z  &       ;Z  &       ;Z  &       R�  &       R�  &       R�  &       R�  &       B�  &       B�  &       B�  &       B�  &       �X  &       �X  &       �X  &       �X  &       �X  &       �X  &       �X  &       �X  &       �0  &       �0  &       �0  &       �0                                                  &       ��  &       ��  &       ��  &       ��  &       �  &       �  &       �  &       �  &       0S &       0S &       0S &       0S &       0S &       0S &       0S &       0S                                                 &       �  &       �  &       �  &       �  &       �:  &       �:  &       �:  &       �:                                                  &       D- &       D- &       D- &       D- &       2�  &       2�  &       2�  &       2�  &       Z  &       Z  &       Z  &       Z  &       b:  &       b:  &       b:  &       b:  &       ��  &       ��  &       ��  &       ��  &       �  &       �  &       �  &       �  &       b�  &       b�  &       b�  &       b�  &       D- &       D- &       D- &       D- &       2�  &       2�  &       2�  &       2�  &       #Y  &       #Y  &       #Y  &       #Y                                                                                                  &       �  &       �  &       �  &       �                                                  &       �#  &       �#  &       �#  &       �#  &       �  &       �  &       �  &       �  &       �#  &       �#  &       �#  &       �#  &       ��  &       ��  &       ��  &       ��  &       �  &       �  &       �  &       �  &       ��  &       ��  &       ��  &       ��                                                                                                  &       �  &       �  &       �  &       �  &       Ҩ  &       Ҩ  &       Ҩ  &       Ҩ  &       �  &       �  &       �  &       �  &       >�  &       >�  &       >�  &       >�  &       �  &       �  &       �  &       �  &       Ũ  &       Ũ  &       Ũ  &       Ũ  &       Ũ  &       Ũ  &       Ũ  &       Ũ  &       ��  &       ��  &       ��  &       ��  &       c &       c &       c &       c &       c &       c &       c &       c &       c &       c &       c &       c &       c &       c &       c &       c &       �d &       �d &       �d &       �d                                                                                                                                                 &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �#  &       �#  &       �#  &       �#                                                                                                  &       �#  &       �#  &       �#  &       �#  &       �c &       �c &       �c &       �c &       c &       c &       c &       c &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       n�  &       n�  &       n�  &       n�                                                                                                  &       ��  &       ��  &       ��  &       ��  &       qd &       qd &       qd &       qd &       s%  &       s%  &       s%  &       s%  &       �  &       �  &       �  &       �  &       �#  &       �#  &       �#  &       �#  &       Vc &       Vc &       Vc &       Vc &       c &       c &       c &       c &       ��  &       ��  &       ��  &       ��                                                  &       �#  &       �#  &       �#  &       �#  &       �  &       �  &       �  &       �  &       ~$  &       ~$  &       ~$  &       ~$                                                  &       c &       c &       c &       c &       �  &       �  &       �  &       �  &       �#  &       �#  &       �#  &       �#  &       c &       c &       c &       c &       �#  &       �#  &       �#  &       �#                                                  &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �%                                                                                                                                                 &       �% &       �% &       �% &       �%                                                                                                 &       F& &       F& &       F& &       F& &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �%                                                                                                 &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       E& &       E& &       F& &       F& &       �% &       �% &       �% &       �% &       F& &       F& &       F& &       F& &       �' &       �' &       �' &       �'                                                 &       �% &       �% &       �% &       �% &       F& &       F& &       F& &       F&                                                                                                                                                                                                 &       �% &       �% &       �% &       �%                                                 &       �' &       �' &       �' &       �' &       F& &       F& &       F& &       F& &       �% &       �% &       �% &       �%                                                 &       �% &       �% &       �% &       �% &       F& &       F& &       F& &       F& &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �' &       �' &       �' &       �' &       F& &       F& &       F& &       F&                                                                                                                                                 &       �% &       �% &       �% &       �%                                                 &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �%                                                 &       �% &       �% &       �% &       �%                                                 &       �% &       �% &       �% &       �% &       E& &       E& &       E& &       E& &       F& &       F& &       F& &       F& &       E& &       E& &       E& &       E& &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �% &       �%                                                                                                                                                 &       E& &       E& &       E& &       E&                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �6  &       �6  &       �6  &       �6                                                                                                  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A                                                  &       �6  &       �6  &       �6  &       �6  &       �  &       �  &       �  &       �                                                                                                                                                  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A                                                                                                  &       �6  &       �6  &       �6  &       �6  &       �  &       �  &       �  &       �                                                  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A                                                                                                                                                                                                  &       �  &       �  &       �  &       �  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A                                                                                                                                                  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A  &       �A                                                                                                                                                                                                  &       �A  &       �A  &       �A  &       �A  &       �  &       �  &       �  &       �                                                                                                                                                                                                                                                                                                  &       �A  &       �A  &       �A  &       �A                                                                                                  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �                                                                                                                                                                                                  &       B  &       B  &       B  &       B  &       �  &       �  &       �  &       �  &       J  &       J  &       J  &       J  &       ��  &       ��  &       ��  &       ��  &       �  &       �  &       �  &       �  &       �2  &       �2  &       �2  &       �2                                                  &       �2  &       �2  &       �2  &       �2  &       w  &       w  &       w  &       w  &       B  &       B  &       B  &       B  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       B  &       B  &       B  &       B  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �  &       �  &       �  &       �  &       B  &       B  &       B  &       B                                                  &       ��  &       ��  &       ��  &       ��  &       �  &       �  &       �  &       �  &       w  &       w  &       w  &       w  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       B  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       ��  &       ��  &       ��  &       ��  &       w  &       w  &       w  &       w                                                  &       J  &       J  &       J  &       J                                                                                                                                                                                                  &       �  &       �  &       �  &       �                                                  &       � &       � &       � &       � &       � &       � &       � &       � &       Z�  &       Z�  &       Z�  &       Z�  &       � &       � &       � &       �                                                                                                 &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       +i  &       +i  &       +i  &       +i  &       +i  &       +i  &       +i  &       +i  &       �x  &       �x  &       �x  &       �x  &        &        &        &                                                        &       �I  &       �I  &       �I  &       �I  &       z�  &       z�  &       z�  &       z�  &       +i  &       +i  &       +i  &       +i  &       xx  &       xx  &       xx  &       xx  &       xx  &       xx  &       xx  &       xx  &       �2  &       �2  &       �2  &       �2  &       B  &       B  &       B  &       B  &       w  &       w  &       w  &       w  &       �  &       �  &       �  &       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       r  &       r  &       r  &       r  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �                                                                                                                                                  &       �  &       �  &       �  &       �  &       2  &       2  &       2  &       2  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �                                                                                                  &       �  &       �  &       �  &       �                                                                                                                                                                                                                                                                                                                                                  &       �  &       �  &       �  &       �  &       R  &       R  &       R  &       R  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �                                                  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �                                                  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       2  &       2  &       2  &       2  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �                                                                                                  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �                                                  &       �  &       �  &       �  &       �  &       R  &       R  &       R  &       R  &       b  &       b  &       b  &       b  &       R  &       R  &       R  &       R                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  &       ^�  &       ^�  &       ^�  &       ^�                                                  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D                                                                                                  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       ^�  &       ^�  &       ^�  &       ^�                                                  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D                                                  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       ]�  &       ]�  &       ]�  &       ]�  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D                                                  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D                                                                                                                                                                                                                                                                                                  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D                                                  &       ]�  &       ]�  &       ]�  &       ]�                                                  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�                                                                                                  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�                                                  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       ]�  &       �D  &       �D  &       �D  &       �D                                                                                                                                                                                                  &       �D  &       �D  &       �D  &       �D                                                  &       �D  &       �D  &       �D  &       �D                                                                                                                                                                                                                                                  &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       <  &       <  &       <  &       <  &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       <  &       <  &       <  &       <  &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       <  &       <  &       <  &       <  &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       >  &       >  &       >  &       >  &       ?  &       ?  &       ?  &       ?  &       A  &       A  &       A  &       A  &       B  &       B  &       B  &       B                                                  &       =  &       =  &       =  &       =  &       ?  &       ?  &       ?  &       ?  &       @  &       @  &       @  &       @  &       <  &       <  &       <  &       <  &       =  &       =  &       =  &       =  &       >  &       >  &       >  &       >  &       ?  &       ?  &       ?  &       ?  &       @  &       @  &       @  &       @  &       <  &       <  &       <  &       <  &       =  &       =  &       =  &       =  &       �   &       �   &       �   &       �   &       F  &       F  &       F  &       F  &       =  &       =  &       =  &       =  &       >  &       >  &       >  &       >  &       ?  &       ?  &       ?  &       ?  &       @  &       @  &       @  &       @  &       <  &       <  &       <  &       <  &       =  &       =  &       =  &       =  &       F  &       F  &       F  &       F  &       <  &       <  &       <  &       <  &       =  &       =  &       =  &       =  &       >  &       >  &       >  &       >  &       ?  &       ?  &       ?  &       ?  &       @  &       @  &       @  &       @  &       =  &       =  &       =  &       =  &       F  &       F  &       F  &       F                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       :  &       :  &       :  &       :  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       :  &       :  &       :  &       :  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9                                                  &       9  &       9  &       9  &       9                                                                                                                                                  &       9  &       9  &       9  &       9                                                  &       9  &       9  &       9  &       9                                                  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9                                                  &       9  &       9  &       9  &       9                                                  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9                                                  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9  &       9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  &       �#  &       �#  &       �#  &       �#                                                  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                                                                                                                                                                  &       �#  &       �#  &       �#  &       �#                                                  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                                                                  &       �#  &       �#  &       �#  &       �#                                                                                                  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                                                                                                                  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                                                                                                                                                                                                                  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                                                                                                                  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                                                                                                                  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                                                                  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#  &       �#                                                                                                     b@ �.     b@ �.    �@ A    �@ A    A �I    A �I    �@ �    �@ �    �@ R�    �@ R�                            �@ �     �@ �     "A �D    "A �D                            �A �    �A �                                                                            �s ;    �s ;    �s �^    �s �^                            t �    t �                                                                            _t �    _t �                            �t Ѡ    �t Ѡ                            �t Di    �t Di                            �t �k    �t �k    �t 5	    �t 5	    "u ��    "u ��    �u �    �u �    �u =    �u =    "v �    "v �    Bv �    Bv �    Mv �    Mv �    bv d    bv d                                                    �w ^    �w ^                            �w Dq    �w Dq                                                                            �x     �x     =y �    =y �    �y �    �y �    �y ��    �y ��    �y �%    �y �%    �v D    �v D  "       m  "       m  "  �A m  "  �A m  "       m  "       m  "       m  "       m  "       m  "       m  "  �B m  "  �B m  "       m  "       m  "       m  "       m  "       m  "       m  "  eC m  "  eC m  "       m  "       m  "       m  "       m  "       m  "       m  "  �E m  "  �E m  "       m  "       m  "       m  "       m  "       �  "       �  "  �F �  "  �F �  "       �  "       �  "       �  "       �  "       �  "       �  "  �G �  "  �G �  "       �  "       �  "       �  "       �  "       �  "       �  "  �I �  "  �I �  "       �  "       �  "       �  "       �  "       �  "       �  "  L �  "  L �  "       �  "       �  "       �  "       �  "       A  "       A  "  �Q A  "  �Q A  "       A  "       A  "       A  "       A  "       A  "       A  "  �R A  "  �R A  "       A  "       A  "       A  "       A  "       A  "       A  "  ES A  "  ES A  "       A  "       A  "       A  "       A  "       A  "       A  "  �U A  "  �U A  "       A  "       A  "       A  "       A  "       �   "       �   "  �N �   "  �N �   "       �   "       �   "       �   "       �   "       �   "       �   "  O �   "  O �   "       �   "       �   "       �   "       �   "       �   "       �   "  �O �   "  �O �   "       �   "       �   "       �   "       �   "       �   "       �   "  �P �   "  �P �   "       �   "       �   "       �   "       �   "       R�  "       R�  "  �W R�  "  �W R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "  Y R�  "  Y R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "  Z R�  "  Z R�  "       R�  "       R�  "       R�  "       R�  "       R�  "       R�  "  ,[ R�  "  ,[ R�  "       R�  "       R�  "       R�  "       R�  "       �I  "       �I  "  �\ �I  "  �\ �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "  Y] �I  "  Y] �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "  @_ �I  "  @_ �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "  �` �I  "  �` �I  "       �I  "       �I  "       �I  "       �I  "       �D  "       �D  "  |b �D  "  |b �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "  {c �D  "  {c �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "  �d �D  "  �d �D  "       �D  "       �D  "       �D  "       �D  "       �D  "       �D  "  #g �D  "  #g �D  "       �D  "       �D  "       �D  "       �D                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       �  "       �  "  �p �  "  �p �  "       �  "       �  "       �  "       �  "       �  "       �  "  Nq �  "  Nq �  "       �  "       �  "       �  "       �  "       �  "       �  "  )r �  "  )r �  "       �  "       �  "       �  "       �  "       �  "       �  "  �r �  "  �r �  "       �  "       �  "       �  "       �  "       s  "       s  "       s  "       s  "       s  "       s  "       s  "       s  "       �  "       �  "         "         "         "         "         "         "       '  "       '  "       o  "       o  "       �  "       �  "       �  "       �  "       #  "       #  "       G  "       G  "       k  "       k  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       N	  "       ~	  "       ~	  "       ~	  "       ~	  "       ~	  "       ~	  "       ~	  "       ~	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       
  "       
  "       
  "       
  "       
  "       
  "       &
  "       &
  "       2
  "       2
  "       >
  "       >
  "       J
  "       J
  "       b
  "       b
  "       n
  "       n
  "       z
  "       z
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       
  "       
  "         "         "       "  "       "  "       .  "       .  "       :  "       :  "       F  "       F  "       R  "       R  "       ^  "       ^  "       j  "       j  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "       +  "       +  "       7  "       7  "       C  "       C  "       O  "       O  "       [  "       [  "       g  "       g  "       s  "       s  "         "         "       �  "       s  "       s  "       s  "       s  "       s  "       s  "       s  "       s  "       s  "       s  "       s  "       �  "       CB  "         "         "       '  "       �B  "       o  "       o  "       �  "       �  "       �  "       cC  "       #  "       �C  "       G  "       �C  "       k  "       �C  "       �  "       ob  "       �  "       ;D  "       �  "       �  "       _  "       �  "       `  "       �  "       a  "       �  "       b  "       �  "       c  "       �  "       �  "       �  "       e  "       �  "       f  "       �  "       g  "       �  "       h  "       �  "       i  "       �  "       j  "       �  "       �  "       �  "       �  "       k  "       N	  "       ~	  "       ~	  "       ~	  "       ~	  "       ~	  "       ~	  "       ~	  "       ~	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       
  "       
  "       
  "       �  "       
  "       
  "       &
  "       &
  "       2
  "       2
  "       >
  "       >
  "       J
  "       J
  "       b
  "       �  "       n
  "       n
  "       z
  "       z
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       ?  "       �
  "       K  "       �
  "       W  "       �
  "       c  "       �
  "          "       
  "       �  "         "       �  "       "  "       �  "       .  "       �  "       :  "         "       F  "       F  "       R  "       R  "       ^  "       ^  "       j  "       j  "       v  "       v  "       �  "         "       �  "         "       �  "       t  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       G  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       w  "         "       �  "         "       �  "         "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "       +  "       +  "       7  "       �  "       C  "       C  "       O  "       O  "       [  "       [  "       g  "       �  "       s  "       �  "         "       �  "       �  "       s  "       s  "       y  "       y  "         "         "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "       	  "       	  "         "         "         "         "         "         "       !  "       !  "       '  "       '  "       -  "       -  "       3  "       3  "       9  "       9  "       ?  "       ?  "       E  "       E  "       K  "       K  "       Q  "       Q  "       W  "       W  "       ]  "       ]  "       c  "       c  "       i  "       i  "       o  "       o  "       u  "       u  "       {  "       {  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "         "         "         "         "       #  "       #  "       )  "       )  "       /  "       /  "       5  "       5  "       ;  "       ;  "       A  "       A  "       G  "       G  "       M  "       M  "       S  "       S  "       Y  "       Y  "       _  "       _  "       e  "       e  "       k  "       k  "       q  "       q  "       w  "       w  "       }  "       }  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       v  "       v  "       |  "       |  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "        	  "        	  "       	  "       	  "       	  "       	  "       	  "       	  "       	  "       	  "       	  "       	  "       $	  "       $	  "       *	  "       *	  "       0	  "       0	  "       6	  "       6	  "       <	  "       <	  "       B	  "       B	  "       H	  "       H	  "       N	  "       N	  "       T	  "       T	  "       Z	  "       Z	  "       `	  "       `	  "       f	  "       f	  "       l	  "       l	  "       r	  "       r	  "       x	  "       x	  "       ~	  "       ~	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       
  "       
  "       
  "       
  "       
  "       
  "       
  "       
  "       
  "       
  "        
  "        
  "       &
  "       &
  "       ,
  "       ,
  "       2
  "       2
  "       8
  "       8
  "       >
  "       >
  "       D
  "       D
  "       J
  "       J
  "       P
  "       P
  "       V
  "       V
  "       \
  "       \
  "       b
  "       b
  "       h
  "       h
  "       n
  "       n
  "       t
  "       t
  "       z
  "       z
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "         "         "       
  "       
  "         "         "         "         "         "         "       "  "       "  "       (  "       (  "       .  "       .  "       4  "       4  "       :  "       :  "       @  "       @  "       F  "       F  "       L  "       L  "       R  "       R  "       X  "       X  "       ^  "       ^  "       d  "       d  "       j  "       j  "       p  "       p  "       v  "       v  "       |  "       |  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "          "          "         "         "         "         "         "         "         "         "         "         "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "         "         "         "         "         "         "       %  "       %  "       +  "       +  "       1  "       1  "       7  "       7  "       =  "       =  "       C  "       C  "       I  "       I  "       O  "       O  "       U  "       U  "       [  "       [  "       a  "       a  "       g  "       g  "       m  "       m  "       s  "       s  "       y  "       y  "         "         "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       s  "       s  "       s  "       s  "       s  "       s  "       s  "         "       �  "       �  "       �  "       �  "       �  "       �  "         "         "       '  "       3  "       K  "       W  "       o  "       o  "       o  "       o  "       o  "       o  "       o  "       {  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "       #  "       /  "       G  "       S  "       k  "       w  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       	  "       	  "       6	  "       B	  "       Z	  "       Z	  "       Z	  "       Z	  "       Z	  "       Z	  "       Z	  "       f	  "       ~	  "       ~	  "       ~	  "       ~	  "       ~	  "       ~	  "       ~	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       �	  "       
  "       
  "       2
  "       >
  "       V
  "       b
  "       z
  "       z
  "       z
  "       z
  "       z
  "       z
  "       z
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       �
  "       
  "         "       .  "       :  "       R  "       ^  "       v  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "       �  "       �  "       �  "       �  "       �  "       �  "         "         "       7  "       7  "       7  "       7  "       7  "       7  "       7  "       C  "       [  "       [  "       [  "       [  "       [  "       [  "       [  "       g  "         "         "         "         "         "         "         "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "       ,  "       2  "       2  "       2  "       2  "       2  "       2  "       2  "       2  "       3  "       3  "       4  "       4  "       5  "       5  "       6  "       7  "       8  "       8  "       9  "       9  "       :  "       :  "       ;  "       ;  "       <  "       =  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       D  "       J  "       J  "       P  "       V  "       V  "       b  "       b  "       h  "       h  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "       "  "       "  "       .  "       .  "       @  "       @  "       R  "       R  "       R  "       R  "       R  "       R  "       R  "       R  "       S  "       S  "       T  "       T  "       U  "       U  "       V  "       W  "       X  "       X  "       Y  "       Y  "       Z  "       Z  "       [  "       [  "       \  "       ]  "       ^  "       ^  "       ^  "       ^  "       ^  "       ^  "       ^  "       ^  "       p  "       p  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "          "          "         "         "         "         "         "         "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "       �#  "         "         "         "         "       �#  "         "       �#  "          "       �#  "       &  "       ,  "       ,  "       2  "       2  "       8  "       8  "       >  "       $  "       D  "       J  "       $  "       P  "       V  "       V  "       \  "       b  "       '$  "       h  "       -$  "       n  "       t  "       9$  "       z  "       ?$  "       �  "       E$  "       �  "       �  "       �  "       �  "       W$  "       �  "       ]$  "       �  "       c$  "       �  "       u$  "       �  "       �$  "       �  "       U;  "       �  "       ��  "       �  "       �  "       �  "       �  "         "         "       "  "       �$  "       .  "       �$  "       @  "       @  "       X  "       ^  "       ^  "       ^  "       ^  "       #%  "       p  "       p  "       �  "       �  "       �  "       S%  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "          "          "         "         "         "         "         "         "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "         "         "         "          "          "       &  "       ,  "       ,  "       2  "       2  "       8  "       8  "       >  "       >  "       D  "       J  "       J  "       P  "       V  "       V  "       \  "       b  "       b  "       h  "       h  "       n  "       t  "       t  "       z  "       z  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "       
  "       
  "         "         "         "         "         "       "  "       (  "       .  "       .  "       4  "       :  "       :  "       @  "       F  "       F  "       L  "       L  "       R  "       X  "       ^  "       ^  "       d  "       j  "       j  "       p  "       v  "       v  "       |  "       |  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "          "         "         "         "         "         "         "         "         "         "         "       $  "       *  "       *  "       0  "       0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "          "       &  "       ,  "       ,  "       ,  "       ,  "       2  "       8  "       >  "       >  "       >  "       >  "       D  "       J  "       P  "       V  "       \  "       b  "       h  "       n  "       t  "       z  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "       
  "         "         "         "         "         "         "         "         "         "       "  "       (  "       .  "       4  "       :  "       @  "       F  "       F  "       F  "       F  "       L  "       L  "       L  "       L  "       R  "       R  "       R  "       R  "       X  "       X  "       X  "       X  "       ^  "       ^  "       ^  "       ^  "       d  "       j  "       p  "       v  "       v  "       v  "       v  "       |  "       |  "       |  "       |  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "          "         "         "         "         "         "         "         "         "       $  "       *  "       0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "         "         "         "         "         "         "       O  "       U  "       U  "       g  "       m  "       m  "         "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "       '  "       -  "       -  "       ?  "       E  "       E  "       Q  "       ]  "       ]  "       i  "       o  "       o  "       {  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "         "         "         "         "         "         "       O  "       U  "       U  "       g  "       m  "       m  "         "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "       '  "       -  "       -  "       ?  "       E  "       E  "       Q  "       ]  "       ]  "       i  "       o              "       {  "       �              "       �              "       �              "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "         "         "         "         "         "         "       %  "       %  "       1  "       1  "       =  "       =  "       I  "       I  "       U  "       a  "       a  "       m  "       m  "       y  "       y  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       	  "       	  "         "       !  "       !  "       -  "       -  "       9  "       9  "       E  "       E  "       Q  "       Q  "       ]  "       ]  "       i  "       i  "       u  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "         "         "         "         "         "         "         "         "         "       %  "       1  "       =  "       =  "       =  "       =  "       I  "       I  "       I  "       I  "       U  "       a  "       m  "       m  "       m  "       m  "       y  "       y  "       y  "       y  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       	  "       	  "       	  "       	  "         "       !  "       -  "       -  "       -  "       -  "       9  "       9  "       9  "       9  "       E  "       E  "       E  "       E  "       Q  "       ]  "       ]  "       ]  "       ]  "       i  "       i  "       i  "       i  "       u  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "         "         "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       k  "       k  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "       h  "       h  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "       (  "       (  "       L  "       L  "       p  "       p  "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       k  "       k  "       k  "       k  "       ��  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "       h  "       *  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "       �R  "       (  "       -  "       L  "       L  "       p  "       p  "       �  "       M                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "       G  "       G  "       M  "       S  "       S  "       Y  "       _  "       _  "       e  "       k  "       k  "       q  "       w  "       w  "       }  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "         "          "          "       &  "       ,  "       ,  "       2  "       8  "       8  "       >  "       D  "       D  "       J  "       P  "       P  "       V  "       \  "       \  "       b  "       h  "       h  "       n  "       t  "       t  "       z  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "       
  "         "         "         "         "         "       "  "       (  "       (  "       .  "       4  "       4  "       :  "       @  "       @  "       F  "       L  "       L  "       R  "       X  "       X  "       ^  "       d  "       d  "       j  "       p  "       p  "       v  "       |  "       |  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       G  "       G  "       G  "       G  "       G  "       G  "       G  "       S  "       _  "       _  "       _  "       _  "       k  "       k  "       k  "       k  "       w  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "          "          "          "          "       ,  "       ,  "       ,  "       ,  "       8  "       D  "       P  "       P  "       P  "       P  "       \  "       \  "       \  "       \  "       h  "       t  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "         "         "         "       (  "       4  "       @  "       @  "       @  "       @  "       L  "       L  "       L  "       L  "       X  "       d  "       p  "       p  "       p  "       p  "       |  "       |  "       |  "       |  "       �  "       �  "       �  "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       _�  "       _�  "       g�  "       g�  "       o�  "       o�  "       o�  "       o�  "       o�  "       w�  "       w�  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ǻ  "       ǻ  "       ϻ  "       ϻ  "       ϻ  "       ϻ  "       ϻ  "       ׻  "       ׻  "       ߻  "       ߻  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       '�  "       '�  "       /�  "       /�  "       7�  "       7�  "       ?�  "       ?�  "       G�  "       G�  "       O�  "       O�  "       W�  "       W�  "       _�  "       _�  "       g�  "       g�  "       o�  "       o�  "       w�  "       w�  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       Ǽ  "       Ǽ  "       ϼ  "       ϼ  "       ׼  "       ׼  "       ׼  "       ׼  "       ׼  "       ߼  "       ߼  "       �  "       �  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       '�  "       '�  "       /�  "       /�  "       7�  "       7�  "       ?�  "       ?�  "       G�  "       G�  "       O�  "       O�  "       W�  "       W�  "       _�  "       _�  "       g�  "       g�  "       o�  "       o�  "       w�  "       w�  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       <9  "       <9  "       D9  "       D9  "       L9  "       L9  "       T9  "       T9  "       \9  "       \9  "       d9  "       d9  "       l9  "       l9  "       t9  "       t9  "       |9  "       |9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       :  "       $:  "       $:  "       ,:  "       ,:  "       4:  "       4:  "       <:  "       <:  "       D:  "       D:  "       D:  "       D:  "       D:  "       L:  "       L:  "       T:  "       T:  "       \:  "       \:  "       \:  "       \:  "       \:  "       \:  "       \:  "       \:  "       `:  "       `:  "       d:  "       d:  "       h:  "       h:  "       l:  "       l:  "       p:  "       p:  "       t:  "       t:  "       t:  "       t:  "       t:  "       |:  "       |:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "        ;  "        ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       $;  "       $;  "       ,;  "       ,;  "       ,;  "       ,;  "       ,;  "       4;  "       4;  "       <;  "       D;  "       D;  "       L;  "       T;  "       T;  "       \;  "       \;  "       d;  "       d;  "       d;  "       d;  "       d;  "       l;  "       t;  "       t;  "       |;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       _�  "       _�  "       g�  "       g�  "       o�  "       o�  "       o�  "       o�  "       o�  "       w�  "       w�  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       d�  "       ��  "       ��  "       ��  "       ��  "       l�  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ǻ  "       ǻ  "       ϻ  "       ϻ  "       ϻ  "       ϻ  "       ϻ  "       ׻  "       ׻  "       ߻  "       ߻  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       '�  "       '�  "       /�  "       /�  "       7�  "       7�  "       ?�  "       ?�  "       G�  "       G�  "       O�  "       O�  "       W�  "       W�  "       _�  "       _�  "       g�  "       g�  "       o�  "       o�  "       w�  "       w�  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       Ǽ  "       Ǽ  "       ϼ  "       ϼ  "       ׼  "       ׼  "       ��  "       ��  "       ��  "       ��  "       �  "       �  "       '�  "       ��  "       /�  "       ��  "       7�  "       �  "       W�  "       $�  "       _�  "       ��  "       g�  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       D9  "       %>  "       L9  "       L9  "       T9  "       T9  "       t9  "       t9  "       |9  "       |9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       :  "       :  "       ,:  "       ,:  "       D:  "       D:  "       D:  "       D:  "       D:  "       L:  "       L:  "       T:  "       T:  "       \:  "       \:  "       \:  "       \:  "       \:  "       d:  "       d:  "       l:  "       l:  "       t:  "       t:  "       t:  "       t:  "       t:  "       �:  "       m?  "       �:  "       �:  "       �:  "       �?  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �?  "       �:  "       �?  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �?  "       �:  "       �?  "       ;  "       ;  "       ;  "       ;  "       �?  "       ;  "       ;  "       ;  "       ;  "       $;  "       $I  "       ,;  "       ,;  "       4;  "       4;  "       4;  "       4;  "       4;  "       <;  "       D;  "       D;  "       L;  "       T;  "       T;  "       \;  "       \;  "       d;  "       d;  "       d;  "       d;  "       d;  "       l;  "       t;  "       t;  "       |;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       W�  "       W�  "       _�  "       _�  "       g�  "       g�  "       o�  "       o�  "       w�  "       w�  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ǻ  "       ǻ  "       ϻ  "       ϻ  "       ׻  "       ׻  "       ߻  "       ߻  "       �  "       �  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       '�  "       '�  "       /�  "       /�  "       7�  "       7�  "       ?�  "       ?�  "       G�  "       G�  "       O�  "       O�  "       W�  "       W�  "       _�  "       _�  "       g�  "       g�  "       o�  "       o�  "       w�  "       w�  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       Ǽ  "       Ǽ  "       ϼ  "       ϼ  "       ׼  "       ׼  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       �  "       �  "       �  "       �  "       '�  "       '�  "       +�  "       /�  "       /�  "       3�  "       7�  "       7�  "       G�  "       W�  "       W�  "       [�  "       _�  "       _�  "       c�  "       g�  "       g�  "       w�  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       D9  "       D9  "       H9  "       L9  "       L9  "       P9  "       T9  "       T9  "       d9  "       t9  "       t9  "       x9  "       |9  "       |9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       :  "       :  "       :  "       $:  "       ,:  "       ,:  "       <:  "       D:  "       D:  "       H:  "       L:  "       L:  "       P:  "       T:  "       T:  "       X:  "       \:  "       \:  "       `:  "       d:  "       d:  "       h:  "       l:  "       l:  "       p:  "       t:  "       t:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "        ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       $;  "       $;  "       ,;  "       ,;  "       4;  "       4;  "       <;  "       D;  "       D;  "       L;  "       T;  "       T;  "       \;  "       \;  "       d;  "       d;  "       l;  "       t;  "       t;  "       |;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       W�  "       _�  "       _�  "       _�  "       _�  "       _�  "       _�  "       _�  "       g�  "       o�  "       o�  "       o�  "       o�  "       w�  "       �  "       �  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ǻ  "       ϻ  "       ϻ  "       ϻ  "       ϻ  "       ׻  "       ߻  "       ߻  "       ߻  "       ߻  "       �  "       �  "       �  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       '�  "       /�  "       7�  "       ?�  "       ?�  "       ?�  "       ?�  "       ?�  "       ?�  "       ?�  "       C�  "       G�  "       G�  "       G�  "       G�  "       G�  "       G�  "       G�  "       O�  "       W�  "       _�  "       g�  "       o�  "       o�  "       o�  "       o�  "       o�  "       o�  "       o�  "       s�  "       w�  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ü  "       Ǽ  "       ˼  "       ϼ  "       Ӽ  "       ׼  "       ߼  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       ��  "       ��  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       '�  "       /�  "       7�  "       7�  "       7�  "       7�  "       7�  "       7�  "       7�  "       ?�  "       G�  "       G�  "       G�  "       G�  "       G�  "       G�  "       G�  "       O�  "       W�  "       _�  "       g�  "       g�  "       g�  "       g�  "       g�  "       g�  "       g�  "       o�  "       w�  "       w�  "       w�  "       w�  "       w�  "       w�  "       w�  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       <9  "       D9  "       L9  "       T9  "       T9  "       T9  "       T9  "       T9  "       T9  "       T9  "       \9  "       d9  "       l9  "       t9  "       t9  "       t9  "       t9  "       t9  "       t9  "       t9  "       |9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       �9  "       :  "       :  "       :  "       :  "       $:  "       ,:  "       4:  "       <:  "       D:  "       D:  "       D:  "       D:  "       D:  "       D:  "       D:  "       L:  "       T:  "       \:  "       d:  "       d:  "       d:  "       d:  "       d:  "       d:  "       d:  "       l:  "       l:  "       l:  "       l:  "       l:  "       l:  "       l:  "       p:  "       t:  "       t:  "       t:  "       t:  "       t:  "       t:  "       t:  "       |:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "       �:  "        ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       ;  "       $;  "       ,;  "       4;  "       4;  "       4;  "       4;  "       <;  "       D;  "       L;  "       T;  "       \;  "       d;  "       d;  "       d;  "       d;  "       l;  "       t;  "       |;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �;  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       J  "       J  "       1J  "       1J  "       AJ  "       AJ  "       QJ  "       QJ  "       aJ  "       aJ  "       iJ  "       iJ  "       yJ  "       yJ  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       K  "       K  "       1K  "       1K  "       AK  "       AK  "       QK  "       QK  "       aK  "       aK  "       iK  "       iK  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �X  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       J  "       =Y  "       1J  "       1J  "       AJ  "       AJ  "       QJ  "       QJ  "       aJ  "       aJ  "       iJ  "       iJ  "       yJ  "       yJ  "       yJ  "       yJ  "       yJ  "       {J  "       {J  "       {J  "       {J  "       {J  "       }J  "       }J  "       }J  "       }J  "       }J  "       J  "       J  "       J  "       J  "       J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       ux  "       K  "       K  "       1K  "       1K  "       AK  "       AK  "       QK  "       QK  "       iK  "       iK  "       yK  "       yK  "       yK  "       yK  "       yK  "       {K  "       {K  "       {K  "       {K  "       {K  "       }K  "       }K  "       }K  "       }K  "       }K  "       K  "       K  "       K  "       K  "       K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �i  "       �K  "       �i  "       �K  "       j  "       �K  "       5y  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       �I  "       J  "       	J  "       	J  "       J  "       J  "       J  "       J  "       !J  "       !J  "       )J  "       )J  "       1J  "       9J  "       9J  "       AJ  "       IJ  "       IJ  "       QJ  "       QJ  "       YJ  "       YJ  "       aJ  "       aJ  "       iJ  "       iJ  "       qJ  "       yJ  "       yJ  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       �J  "       K  "       	K  "       	K  "       K  "       K  "       K  "       K  "       !K  "       !K  "       )K  "       )K  "       1K  "       9K  "       9K  "       AK  "       IK  "       IK  "       QK  "       QK  "       YK  "       YK  "       aK  "       aK  "       iK  "       iK  "       qK  "       yK  "       yK  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       �K  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       �I  &       J  &       J  &       J  &       J  &       	J  &       	J  &       	J  &       	J  &       J  &       J  &       !J  &       !J  &       !J  &       !J  &       )J  &       )J  &       )J  &       )J  &       1J  &       9J  &       AJ  &       AJ  &       AJ  &       AJ  &       IJ  &       IJ  &       IJ  &       IJ  &       QJ  &       YJ  &       aJ  &       aJ  &       aJ  &       aJ  &       iJ  &       iJ  &       iJ  &       iJ  &       qJ  &       yJ  &       yJ  &       yJ  &       yJ  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       �J  &       K  &       K  &       K  &       K  &       	K  &       	K  &       	K  &       	K  &       K  &       K  &       !K  &       !K  &       !K  &       !K  &       )K  &       )K  &       )K  &       )K  &       1K  &       9K  &       AK  &       AK  &       AK  &       AK  &       IK  &       IK  &       IK  &       IK  &       QK  &       YK  &       aK  &       aK  &       aK  &       aK  &       iK  &       iK  &       iK  &       iK  &       qK  &       yK  &       yK  &       yK  &       yK  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       �K  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �  &       �  &       ��  &       ��  &       �  &       �  &       �  &       �  &       L�  &       L�  &       ^�  &       ^�  &       |�  &       |�  &       ��  &       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       Ξ  &       Ξ  &       ��  &       ��  &       �  &       �  &       "�  &       "�  &       .�  &       .�  &       ^�  &       2�  &       p�  &       p�  &       ��  &       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      &       �D  &       ��  &       ��  &         &       Ȟ  &       Ȟ  &       Ξ  &       Ԟ  &       Ԟ  &       ��  &       �  &       �  &       �  &       ��  &       ��  &       ��  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       "�  &       (�  &       (�  &       .�  &       4�  &       4�  &       @�  &       F�  &       F�  &       R�  &       X�  &       X�  &       ^�  &       d�  &       d�  &       p�  &       v�  &       v�  &       |�  &       |�  &       ��  &       ��  &       ��  &       ��  &       h�  &       h�  &       t�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       �D  &       Ξ  &       Ԟ  &       Ԟ  &       Ԟ  &       Ԟ  &       ڞ  &       ڞ  &       ڞ  &       ڞ  &       ��  &       �  &       �  &       �  &       ��  &       ��  &       �  &       �  &       �  &       �  &       
�  &       
�  &       
�  &       
�  &       �  &       �  &       �  &       "�  &       (�  &       .�  &       4�  &       4�  &       4�  &       4�  &       :�  &       :�  &       :�  &       :�  &       @�  &       F�  &       L�  &       R�  &       X�  &       ^�  &       d�  &       d�  &       d�  &       d�  &       j�  &       j�  &       j�  &       j�  &       p�  &       v�  &       |�  &       |�  &       |�  &       |�  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       A  &       A  &       Y  &       Y  &       i  &       i  &       y  &       y  &       �  &       �  &       �  &       �  &       I  &       I  &       I  &       I  &       I  &       I  &       I  &       I  &       y  &       y  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       	  &       	  &       9  &       9  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       )  &       )  &       A  &       A  &       Y  &       Y  &       q  &       q  &       �  &       �  &       �  &       �  &       �  &       �  &         &                     &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       �   &       A  &       A  &       Y  &       Y  &       i  &       i  &       y  &       y  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &         &         &         &         &         &         &         &         &         &         &         &         &       %  &       %  &       +  &       +  &       1  &       1  &       7  &       7  &       =  &       =  &       C  &       C  &       I  &       I  &       I  &       I  &       I  &       I  &       I  &       I  &       I  &       I  &       I  &       y  &       y  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       	  &       	  &       9  &       9  &       Q  &       Q  &       i  &       i  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &         &         &       	  &       	  &         &         &         &         &       !  &       !  &       )  &       )  &       1  &       1  &       9  &       9  &       A  &       A  &       I  &       I  &       Q  &       Q  &       Y  &       Y  &       a  &       a  &       i  &       i  &       q  &       q  &       y  &       y  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &         &         &       	  &       	  &         &         &         &         &       !  &       !  &       )  &       )  &       1  &       1  &       7  &       7  &       =  &       =                                      &       �  &       �  &       �  &       �  &       �  &       i   &       i   &       �   &       �   &       )  &       )  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &         &         &         &         &         &         &       %  &       %  &       1  &       1  &       =  &       =  &       I  &       I  &       U  &       U  &       a  &       a  &       m  &       m  &       y  &       y  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       	  &       	  &         &         &       !  &       !  &       -  &       -  &       9  &       9  &       E  &       E  &       Q  &       Q  &       ]  &       ]  &       i  &       i  &       u  &       u  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &         &         &         &         &         &         &       )  &       )  &       5  &       5  &       A  &       A  &       M  &       M  &       Y  &       Y  &       e  &       e  &       q  &       q  &       }  &       }  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &         &         &         &         &         &         &       %  &       %  &       1  &       1  &       =  &       =              &       �  &       i   &       �   &       )  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &         &         &         &         &         &         &         &         &         &         &       %  &       1  &       7  &       =  &       C  &       I  &       I  &       I  &       I  &       I  &       I  &       I  &       U  &       a  &       a  &       a  &       a  &       m  &       m  &       m  &       m  &       y  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       	  &       	  &       	  &       	  &         &       !  &       !  &       !  &       !  &       -  &       -  &       -  &       -  &       9  &       E  &       Q  &       Q  &       Q  &       Q  &       ]  &       ]  &       ]  &       ]  &       i  &       u  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &         &         &         &         &         &         &         &         &         &       )  &       5  &       A  &       A  &       A  &       A  &       M  &       M  &       M  &       M  &       Y  &       e  &       q  &       q  &       q  &       q  &       }  &       }  &       }  &       }  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &         &         &         &         &         &         &         &         &         &       %  &       1  &       1  &       1  &       1  &       =  &       =  &       =  &       =                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          &       ;  &       ;  &       ;  &       ;  &       ;  &       ;  &       ;  &       ;  &       <  &       <  &       =  &       =  &       >  &       >  &       ?  &       ?  &       @  &       @  &       A  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^  &       �^                                                                                                                                                                                                                                                                                      &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �                                                                                                                                                                                                                                                                                                                                                                                                              &       Ѡ  &       Ѡ  &       Ѡ  &       Ѡ  &       Ѡ  &       Ѡ  &       Ѡ  &       Ѡ  &       Ҡ                                                                                                                                      &       Di  &       Di  &       Di  &       Di  &       Di  &       Di  &       Di  &       Di  &       Ei  &       Ei  &       Fi  &       Fi  &       Gi  &       Gi  &       Hi  &       Hi  &       Ii  &       Ii  &       Ji  &       Ji  &       Ki  &       Ki  &       Li  &       Li  &       Mi  &       Mi  &       Ni                                                                                                                                                                                                                                                                                      &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       �k  &       5	  &       5	  &       5	  &       5	  &       5	  &       5	  &       5	  &       5	  &       6	  &       6	  &       7	  &       7	  &       8	  &       8	  &       9	  &       9	  &       :	  &       :	  &       ;	  &       ;	  &       <	  &       <	  &       =	  &       =	  &       >	  &       >	  &       ?	  &       ?	  &       @	  &       @	  &       @	  &       @	  &       @	  &       A	  &       A	  &       B	  &       B	  &       C	  &       C	  &       D	  &       D	  &       E	  &       E	  &       F	  &       F	  &       G	  &       G	  &       H	  &       H	  &       I	  &       I	  &       J	  &       J	  &       K	  &       K	  &       L	  &       L	  &       M	  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ¢  &       ¢  &       â  &       â  &       Ģ  &       Ģ  &       Ţ  &       Ţ  &       Ţ  &       Ţ  &       Ţ  &       Ƣ  &       Ƣ  &       Ǣ  &       Ǣ  &       Ȣ  &       Ȣ  &       ɢ  &       ɢ  &       ɢ  &       ɢ  &       ɢ  &       ʢ  &       ʢ  &       ˢ  &       ˢ  &       ̢  &       ̢  &       ͢  &       ͢  &       ͢  &       ͢  &       ͢  &       ΢  &       ΢  &       Ϣ  &       Ϣ  &       Т  &       Т  &       Ѣ  &       Ѣ  &       Ѣ  &       Ѣ  &       Ѣ  &       Ң  &       Ң  &       Ӣ  &       Ӣ  &       Ԣ  &       Ԣ  &       բ  &       բ  &       բ  &       բ  &       բ  &       ֢  &       ֢  &       ע  &       ע  &       آ  &       آ  &       ڢ  &       ڢ  &       ڢ  &       ڢ  &       ڢ  &       ۢ  &       ۢ  &       ܢ  &       ܢ  &       ݢ  &       ݢ  &       ޢ  &       ޢ  &       ޢ  &       ޢ  &       ޢ  &       ߢ  &       ߢ  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       =  &       =  &       =  &       =  &       =  &       =  &       =  &       =  &       >  &       >  &       j  &       j  &       k  &       k  &       l  &       l  &       l  &       l  &       l  &       n  &       n  &       n  &       n  &       n  &       p  &       p  &       r  &       r  &       t  &       t  &       v  &       v  &       x  &       x  &       z  &       z  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &         &         &         &         &         &         &         &       
  &       
  &         &         &         &         &         &         &          &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �              &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       d  &       d  &       d  &       d  &       d  &       d  &       d  &       d  &       e  &       e  &       f  &       f  &       g  &       g  &       h  &       h  &       i  &       i  &       j  &       j  &       k  &       k  &       l  &       l  &       m  &       m  &       n  &       n  &       o  &       o  &       p  &       p  &       q  &       q  &       r  &       r  &       s  &       s  &       t  &       t  &       t  &       t  &       t  &       u  &       u  &       v  &       v  &       w  &       w  &       x  &       x  &       y  &       y  &       z  &       z  &       {  &       {  &       |  &       |  &       }  &       }  &       ~  &       ~  &         &         &         &         &         &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       D  &       D  &       D  &       D  &       D  &       D  &       D  &       D  &       D  &       D  &       D  &       D  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &        �  &        �  &        �  &        �  &        �  &       !�  &       !�  &       "�  &       "�  &       ^�  &       ^�  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��                                                                                                                                                                                                                                                                                      &       ^  &       ^  &       ^  &       ^  &       ^  &       ^  &       ^  &       ^  &       `  &       `  &       b  &       b  &       d  &       d  &       f  &       f  &       f  &       f  &       f  &       h  &       h  &       j  &       j  &       l  &       l  &       n                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      &       Dq  &       Dq  &       Dq  &       Dq  &       Dq  &       Dq  &       Dq  &       Dq  &       Fq  &       Fq  &       Hq  &       Hq  &       Jq  &       Jq  &       Lq  &       Lq  &       Nq  &       Nq  &       Pq  &       Pq  &       Rq  &       Rq  &       Tq  &       Tq  &       Vq  &       Vq  &       Xq  &       Xq  &       Zq  &       Zq  &       \q  &       \q  &       ^q  &       ^q  &       `q  &       `q  &       bq  &       bq  &       dq                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &         &          &          &       !  &       !  &       "  &       "  &       #  &       #  &       #  &       #  &       #  &       $  &       $  &       %  &       %  &       &  &       &  &       '  &       '  &       '  &       '  &       '  &       (  &       (  &       )  &       )  &       *  &       *  &       +  &       +  &       +  &       +  &       +  &       ,  &       ,  &       -  &       -  &       .  &       .  &       /  &       /  &       0  &       0  &       1  &       1  &       2  &       2  &       3  &       3  &       4  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       z  &       z  &       {  &       {  &       |  &       |  &       |  &       |  &       |  &       }  &       }  &       ~  &       ~  &         &         &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       �  &       :  &       :  &       ;  &       ;  &       ;  &       ;  &       ;  &       <  &       <  &       =  &       =  &       =  &       =  &       =  &       >  &       >  &       >  &       >  &       >  &       ?  &       ?  &       ?  &       ?  &       ?  &       @  &       @  &       A  &       A  &       B  &       B  &       C  &       C  &       D  &       D  &       E  &       E  &       F  &       F  &       G  &       G  &       H  &       H  &       H  &       H  &       H  &       I  &       I  &       J  &       J  &       K  &       K  &       L  &       L  &       M  &       M  &       N  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��  &       ��                                                                                      &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �%  &       �:  &       �:  &       �:  &       �:  &       z;  &       z;  &       �  &       �  &       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    L� �     L� �     l� 9    l� 9    ��     ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           "       �   "       �   "  [� �   "  [� �   "       �   "       �   "       �   "       �   "       �   "       �   "  5� �   "  5� �   "       �   "       �   "       �   "       �   "       �   "       �   "  � �   "  � �   "       �   "       �   "       �   "       �   "       �   "       �   "  .� �   "  .� �   "       �   "       �   "       �   "       �   "       9  "       9  "  �� 9  "  �� 9  "       9  "       9  "       9  "       9  "       9  "       9  "  �� 9  "  �� 9  "       9  "       9  "       9  "       9  "       9  "       9  "  7� 9  "  7� 9  "       9  "       9  "       9  "       9  "       9  "       9  "  r� 9  "  r� 9  "       9  "       9  "       9  "       9  "         "         "  G�   "  G�   "         "         "         "         "         "         "  ��   "  ��   "         "         "         "         "         "         "  ƕ   "  ƕ   "         "         "         "         "         "         "  G[   "  G[   "         "         "         "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "         "         "         "         "         "       $  "       $  "       ,  "       ,  "       4  "       4  "       <  "       <  "       D  "       D  "       L  "       L  "       T  "       T  "       \  "       \  "       d  "       d  "       l  "       l  "       t  "       t  "       |  "       |  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "       ,  "       ,  "       ,  "       ,  "       ,  "       \  "       \  "       t  "       t  "       �  "       �  "       �  "       �  "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "         "         "         "         "         "       $  "       $  "       ,  "       ,  "       4  "       4  "       <  "       <  "       <  "       <  "       <  "       D  "       D  "       L  "       L  "       T  "       T  "       \  "       \  "       d  "       d  "       l  "       l  "       t              "       |              "       �              "       �              "       �              "       �              "       �              "       �              "       �  "       �  "       �  "       �  "       �  "       �  "       �              "       �              "       �  "       �  "       �              "       �              "       �  "       �  "       �  "       �  "         "         "         "         "       4  "       <              "       l  "       l  "       �              "       �  "       �  "       �  "       �  "       �  "       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       �  "       �  "       �  "       �  "       �  "         "         "       l  "       l  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "         "         "         "         "         "         "         "       $  "       $  "       ,  "       ,  "       4  "       D  "       D  "       L  "       \  "       \  "       d  "       d  "       l  "       l  "       t  "       t  "       |  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �   "       �  "       �  "         "         "         "       T  "       \  "       d  "       l  "       t  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "          "         "         "         "         "         "          "       $  "       (  "       ,  "       4  "       D  "       L  "       \  "       d  "       t  "       |  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "         "                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       ^  "       ^  "       n  "       n  "       �  "       �  "       ��  "       ��  "       ͢  "       ͢                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       V  "       V  "       v  "       v  "       �  "       �  "       �  "       �  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          "       >  "       >  "       ~  "       ~  "       ��  "       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "       >  "       >  "       >  "       >  "       >  "       >  "       >  "       N  "       ^  "       ^  "       ^  "       ^  "       n  "       n  "       n  "       n  "       ~  "       �  "       �  "       �  "       �  "       �  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ��  "       ͢  "       ͢  "       ͢  "       ͢                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              "       #  "       #  "       #  "       #  "       #  "       #  "       #  "       #  "       )  "       )  "       /  "       /  "       5  "       5  "       ;  "       ;  "       A  "       A  "       G  "       G  "       G  "       G  "       G  "       M  "       M  "       S  "       S  "       Y  "       Y  "       _  "       _  "       e  "       e  "       k  "       k  "       k  "       k  "       k  "       q  "       q  "       w  "       w  "       }  "       }  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                                                                              "       #  "       #  "       #  "       #  "       #  "       #  "       #  "       )  "       )  "       /  "       /  "       5  "       5  "       ;  "       ;  "       A  "       A  "       G  "       G  "       M  "       M  "       M  "       M  "       M  "       S  "       S  "       Y  "       Y  "       _  "       _  "       e  "       e  "       k  "       k  "       q  "       q  "       q  "       q  "       q  "       w  "       w  "       }  "       }  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �  "       �                                                                                                              "       #  "       #  "       k                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          }          �         �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 1� �                               �                    �                    �                    �                    �                    �                    �                               �                    �                    �                               �                    �                    �                    �                    �                    �                    �                    �                               �         �                    �                    �                    �                    �                �� �                           �� �                           u� �                           � �                               �                    �                    �                    �                � �                           H� �                               �                    �                    �                               �                    �                    ]                     ]                 �� }                                �                     �                     �                     �                 C� �                                �                     �                                                                                             �                     �                     �                     �                     �                     �                     �                     �                     �                                �                     �                     �                                �                     �          �                     �                     �                     �                                �                     �                                �                     �                     �                     �                 �� �                                �                     �                 � ,                           �� �                                                                a� ,                           u� @                           �� @                           � @                               @                d� @                               @                    @                d� @                               @                    @                    @                    @                    @                �� @                               A                d� A                               A                    A                    A                    A                    A                d� A                               A         A         A         A         A                    A                T� A                               A                    A                    A                    A                    A                    A                    A                    A                    A                    A         A                    A                    A                    A                    A                    A                    A         A                    A                    A                    A                    A                    M`                    A                    A                    A                    A                d� A                               A         A         A         A                    A         A         A                    A                    A                �� A                               A                    A                    A                    A                    A         A         A         A         A                    A         A                �� A                               A                    A         A         A                    A                    A         A                    A                    A                    A                    A                    A                    A                    A                    A                    A                    A                    A                    A                    A                    A                    A                    A                    A                    A                �� A                           z� B                               B                    B                    B                    B                �� B                           �� C                           �� C                           �� C                           �� C                           �� C                           |� C                           �� C                           4� C                               C                    C                    C                    C                �� C                               ]                    ]                    ]                    ]                    ]                    ]                � ]                           C� ]                               ]                    ]                                                        ]                    ]                    ]                    ]                    ]                    ^                    ^                    ]                    ]                � ]                               ]                    ]                    ]                    ]                    ]                    ]                �� ]                               ]                    ]                    ]                    ]                �� ]                               ]                    ]                    ]                    ]                �� ]                               ]                    ]                    ]                    ]                �� ]                               ]                    ]                    ]                    ]                �� ]                           �� ]                           �� ]                               ]                    ]                    ]                    �                    ]                    ]                    ]                    ]                �� ]                               ^                    ^                !� ^                           a� �                           d� �                               A         m         e�         �         �A     a� �                                �                     �                     �                     �                 �� �                            z� �                            u� �                            1� �                            �� �                            �� �                            �� �                            �� �                                �                     �                     �                     �                     �                     �                 �� �                                �          ]                d� ]                               ]     �� ]                               ]                    ]                d� ]                               ]         ]                    �                    �                    �                    ]         �         �         ]         �         �                � �                               �                               �         �                    �         @                �� @                               @                               @         @                    @         ]                    ]                    ]                    ]                    j                    ]                               ]                               ]                               ]                               ]                               ]                               ]                               ]                               ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             �                    �                    �                               �         �         �         �         �                               �         �                               �                    �                               �         �         �                    �                    �                               �                    �                               �         �                    �                               �                    �         �                               �         �         �                    �                               �                    �         �                               �         �         �                    �                    �                    �         �                               �         �                    �                               �                    �                    �                               �         �                    �                               �                               �                    �         �                               �         �         �                    �                               �                    �         �                               �         �         �                    �                               �                    �                               �                    �                    �                    �                d� �                               �                    �                               �                               �                d� �                               �                    �                               �                               �         �                    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �                �� �                               �                    �         �                    �                    �                    �                    �                               �         �                    �         �                    �         �                    �                               �                    �                    �                    �         �                    �                               �                    �                               �                    �                               �                ɞ �                               �                               �         �                    �                ɟ �                               �                               �         �                    �                ɠ �                               �                               �         �                    �                ɡ �                               �                               �         �                � �                               �                � �                               �                    �         �                    �         �                    �                               �         }                     }                     }                     }                 � }                                }                     }                 ж }                                }                     }                     }                     }                 �� }                                �                     �          �                     �                     �                 i� �                                �          }                                }                     }                     }                                }                     }          }                     }                     }                 � }                                �                     }                                }          }          }                     }          }                 ɢ }                                }                                }          }                     }          @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         @         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �         �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  K          	          	           	          	          	           	          	           	           	          	           	           	          	           	           	          	           	          	           	           	          	           	           	          	           	          	           	           	          	           	           	          	           	          	           	           	          	           	          	           	          	          	           	          	           	           	   �    	           	           	   A�    	           	                                                                                                                                                                          ��    	           	           	          	           	          	           	          	           	          	           	   ��    	           	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	   �� �   	           	           	       �   	           	       �   	           	   +� �   	           	                  �  	           	       �  	                                                                                                                                                                                                                                                                                                                                                                                                                                   	       �  	           	       �  	           	       �  	           	       �  	           	   C� �  	           	           	   +� �  	           	           	       �  	           	       �  	           	   (� �  	           	           	   |� �  	           	           	   �� �  	           	           	   ]� �  	           	           	       �  	   �� �  	           	           	   �� �  	           	           	       �  	       �  	           	       "  	           	       "  	           	       "  	           	       "  	           	   5� �  	           	           	   m� �  	           	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  }              	       }   	           	       �  	           	       �  	           	   �� �  	           	           	   X� �  	           	           	       }   	           	       }   	           	       C  	           	       C  	           	   �� C  	           	           	   X� D  	           	           	       }   	           	       }   	           	   i� }   	           	                  ~   	           	       ~   	           	       �          ]             	       ]  	       ]  	       ]  	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	       ]  	       ]  	       ]  	           	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       p  	           	       p  	           	       p  	           	       p  	           	       p  	       p  	           	       p  	           	       p  	           	       p  	           	       p  	           	       p  	           	   �� p  	           	           	       J  	           	       J  	           	       J  	           	       J  	           	   �� J  	           	           	       {  	           	       {  	           	       {  	           	         	           	         	         	           	         	           	         	           	         	           	         	           	         	           	         	           	   ��   	           	                                                                                      �� p  	           	           	       p  	       p     �� ]  	           	           	       ]  	       ]  	       C  	           	       C  	       C  	       C  	       C  	       C  	           	       C  	       C  	           	       C  	       C  	           	       C  	           	       C  	       C  	           	       C  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	           	       �  	           	           	       �  	       C  	           	       C  	       C  	           	       C  	           	           	       C  	           	           	       C  	           	       C  	       C  	       C  	       C  	       C  	           	       C  	           	       C  	           	       C  	       C  	       C  	       C  	       C  	           	       C  	       C  	           	       C  	           	           	       C  	       C  	           	       C  	           	           	       C  	           	       C  	           	           	       C  	           	           	       C  	           	       C  	           	       C  	           	       C  	           	           	       C  	       C  	       C  	           	           	       C  	       n  	           	           	       n  	       n  	       n  	           	           	       n  	       C  	           	       C  	           	       C  	           	       C  	           	       �   	           	       �   	           	           	       �   	           	           	   o� �   	           	           	       C  	           	           	       C  	           	           	       C  	       C  	       C  	       C  	       C  	       C  	           	       C  	           	           	       C  	       C  	           	       C  	           	           	       C  	           	       C  	           	           	       C  	           	           	       C  	           	       C  	           	           	       C  	           	       C  	           	                  C  	           	       C  	           	       C  	           	       C  	           	       C  	       C  	       C  	       C  	           	       C  	           	           	       C  	       C  	           	       C  	           	           	       C  	       C  	       C  	       C  	           	       C  	           	           	       C  	       C  	           	       C  	           	           	       C  	           	       C  	           	           	       C  	           	           	       C  	           	   �� C  	           	           	       C  	                  C  	           	           	       C  	           	           	       C  	       C  	       C  	           	       C  	       C  	       C  	           	       C  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	   �� ]  	           	           	       ]  	       ]  	       ]  	           	       ]  	           	       ]  	       ]  	       ]  	       ]  	           	       ]  	       ]  	           	       ]  	           	       ]  	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	       ]  	           	       ]  	           	       ]  	       ]  	           	           	       ]  	           	       ]  	           	           	       ]  	           	       ]  	           	       ]  	           	           	       ]  	           	           	       ]  	           	           	       ]  	           	       ]  	           	       ]  	           	           	       ]  	           	           	       ]  	           	       ]  	           	           	   � ]  	           	           	       i  	           	           	       i  	           	           	       i  	           	       i  	           	                  ]  	           	           	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	           	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	       ]  	       ]  	       ]  	           	       ]  	           	       ]  	           	           	       ]  	           	       ]  	           	       `  	           	           	       `  	           	       �  	       �  	           	       �  	           	       �  	           	       �  	           	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	           	       ]  	       ]  	           	       ]  	           	           	       ]  	           	           	       ]  	       ]  	           	       ]  	           	           	       ]  	           	           	       ]  	       ]  	           	       ]  	           	           	       ]  	           	           	       ]  	       �  	           	           	       �  	           	           	       �  	       �  	           	       �  	           	           	       �  	           	       �  	           	           	       �  	       @  	           	   k� @  	           	           	       @  	           	           	       @  	       @  	           	       @  	           	       @  	           	       @  	           	           	       @  	       @  	           	       @         A             	       A  	       A  	           	       A  	           	           	       A  	           	       A  	           	       A  	           	       A  	       A  	           	       A  	           	           	       A  	           	       A  	           	           	       A  	           	       A  	           	           	       A  	           	       A  	           	       A  	           	       A  	           	           	       A  	       A  	           	       A  	       A  	           	       B  	           	       B  	           	       B  	           	           	       B  	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	           	       B  	       B  	           	       B  	       B  	           	       B  	           	       B  	           	       B  	           	           	       B  	       B  	           	       B  	       B  	           	       B  	       B  	           	       B  	           	           	       B  	       �   	           	       �   	           	       �   	       �   	       �   	           	       �   	           	       �   	           	       �   	           	           	       �   	           	       �   	           	       �   	           	           	       �   	           	       �   	       �   	           	       �   	           	       �   	           	   	� �   	           	           	       �   	                  �   	           	           	       �   	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	   5� �   	           	           	       �   	       �   	       �   	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	       4�  	           	       4�  	       4�  	       4�  	           	       4�  	           	       4�  	           	       4�  	           	           	       4�  	           	       4�  	           	       4�  	           	           	       4�  	           	       4�  	       4�  	           	       4�  	           	       4�  	           	   R� 4�  	           	           	       4�  	                  4�  	           	           	       4�  	       4�  	           	   5� 4�  	           	           	       9�  	       9�  	       9�  	       9�  	           	       H�  	       ,  	           	       ,  	       ,  	       ,  	           	       ,  	           	       ,  	           	       ,  	           	           	       ,  	           	       ,  	           	       ,  	           	           	       ,  	           	       ,  	       ,  	           	       ,  	           	       ,  	           	   �� ,  	           	           	       ,  	                  ,  	           	           	       ,  	       ,  	           	   5� ,  	           	           	       1  	       1  	       1  	       1  	           	       @         C             	       C  	           	       C  	           	       C  	           	   �� C  	           	           	       C  	           	       C  	           	    � C  	           	           	   5� C  	           	           	       H  	           	       H  	       H  	           	       H  	           	       H  	           	   i� \  	           	           	       ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	       C  	           	           	       C  	           	       C  	           	       C  	           	           	       C  	           	       C  	       C  	           	       C  	           	       C  	           	   8� C  	           	           	       H  	                  C  	           	           	       C  	       C  	       C  	           	       C  	       g  	       g  	       g  	           	       g  	           	       g  	           	           	       g  	       g  	           	   i� g  	           	           	       h  	           	       h  	           	   5� h  	           	           	   �� i  	           	           	   i� i  	           	           	       j  	           	       j  	           	   5� j  	           	           	       l  	       l  	       l  	       l  	           	       �  	   �� }   	           	           	       }   	           	       }   	           	       }   	           	       }   	           	       }   	           	   �� }   	           	           	       ~   	   �� B  	           	           	       B  	           	       B  	       B  	           	       B  	           	           	       B  	           	       B  	           	       B  	           	       B  	       B  	           	       B  	           	           	       B  	           	       B  	           	           	       B  	           	       B  	           	           	       B  	           	       B  	           	   �� B  	           	           	       B  	           	           	       B  	       B  	       B  	           	       B  	           	       B  	           	           	       B  	           	       B  	           	           	       B  	           	       B  	           	       B  	           	           	       B  	       B  	           	       B  	           	       B  	           	       B  	       B  	           	       B  	       B  	           	       B  	           	           	       B         B             	       B  	           	       B  	           	       B  	           	       B  	           	   T� B  	           	           	   �� B  	           	           	       C  	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	   T� �   	           	           	       �   	           	       �   	       �   	           	       �   	       �   	           	       �   	           	   �� �   	           	           	       �   	       B  	           	       B  	       B  	           	       B  	           	       B  	           	           	       B  	           	       B  	       B  	           	       B  	           	       B  	           	       B  	       B  	           	       B  	           	           	       B  	           	       B  	       B  	           	       B  	       B  	           	       B  	       B  	           	       B  	           	       B  	           	       B  	           	       B  	       B  	       B  	           	       B  	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	           	       B  	           	       B  	           	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	       B  	       B  	       B  	           	       B  	           	           	       B  	       B  	           	       B  	           	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	           	       B  	           	       B  	       B  	           	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	       B  	       B  	       B  	       B  	       B  	           	       B  	           	           	       B  	       B  	           	       B  	           	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       B  	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       B  	           	       C  	       C  	           	       C  	       C  	           	       C  	           	       C  	       C  	           	       C  	           	       C  	           	       C  	           	       C  	       C  	       C  	           	       C  	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	                  C  	           	       C  	           	       C  	           	       C  	       C  	           	       C  	       C  	           	       C  	           	       C  	           	       C  	       C  	           	       C  	       C  	           	       C  	           	       C  	           	       C  	       C  	           	       C  	       C  	           	       C  	           	       C  	           	       C  	       C  	           	       C  	       C  	           	       C  	           	       C  	           	           	       C  	           	       C  	           	           	       C  	           	       C  	           	           	       C  	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	       C  	           	       C  	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	   �� C  	           	           	       C  	       C  	           	       C  	       C  	           	       C  	       C  	           	       C  	           	           	       C  	   �� �I  	           	           	       �I  	           	       �I  	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	       �I  	       �I  	           	       �I  	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	   3� �I  	           	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	   �� :  	           	           	       :  	           	       :  	       :  	           	       :  	           	       :  	           	       :  	           	       :  	       :  	       :  	           	       :  	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	   \� :  	           	           	       ;  	           	       ;  	           	       ;  	           	       ;  	           	       ;  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       ;  	           	       ;  	           	       ;  	           	       J  	   �� �  	           	           	       �  	           	       �  	           	       �  	           	       �  	       �  	           	       �  	           	   � �  	           	           	         	           	         	                  �  	           	       �  	       �  	           	       �  	           	       �  	           	       �  	           	       �  	       �  	       �  	           	       �  	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	   3� �  	           	           	       �  	       �  	           	       �  	       �  	           	       �  	           	    �  �  	           	           	       �  	           	       �  	           	   �  �  	           	           	       �  	           	       �  	           	   T� �  	           	           	   q� �  	           	           	       �  	           	       �  	           	    �  �  	           	           	       �  	       �  	           	   �  �  	           	           	       �  	       :  	           	       :  	           	   T� :  	           	           	       :  	           	       :  	       :  	           	       :  	       :  	           	       :  	           	   q� :  	           	           	       ;  	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	       �  	       �  	       �  	           	       �  	           	           	       �  	       �  	           	       �  	           	           	       �  	       �  	           	       �  	           	           	       �  	       �  	           	       �  	           	           	       �  	           	       �  	       �  	       �  	           	       �  	           	       �  	       �  	           	       �  	           	       �  	           	       �  	       �  	       �  	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	           	       �  	       �  	           	       �  	           	       �  	           	       �  	       �  	           	       �  	       �  	       �  	       �  	       �  	           	           	       �  	           	       �  	       �  	           	       �  	           	           	       �  	           	           	       �  	           	       �  	           	       �  	           	       �  	           	           	       �  	           	           	       �  	       �  	       �  	           	       �  	           	   �� �  	           	           	       �     �� @                        	   �� A  	           	           	   	� A  	           	           	   �� A  	           	           	       A  	   �� �   	           	           	   	� �   	           	           	   �� �   	           	           	       �   	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	           	       A  	           	   � A  	           	           	       A  	           	       A  	           	       A  	           	       A  	           	           	       A  	           	       A  	           	       A  	           	           	       A  	       A  	           	       A  	           	           	       A  	           	       A  	           	           	       A  	       A  	           	       A  	           	           	       A  	       A  	           	       A  	           	       A  	           	       I 	           	       I 	           	           	       I 	           	   p� I 	           	           	       A  	                  A  	           	           	       A  	           	       A  	           	       A  	           	       �  	           	       �  	       �  	       �  	       �  	           	       �  	           	       �  	           	       �  	           	       A  	           	       A  	           	   .� A  	           	           	       A  	           	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	           	       A  	       A  	           	       A  	           	       A  	           	       A  	           	           	       A  	       A  	           	       A  	           	       A  	           	       A  	           	           	       A  	       A  	           	       A  	           	       A  	       @  	           	       @  	       @  	           	       @  	           	       @  	           	       @  	           	   �� @  	           	           	       A  	           	       A  	           	       A  	       A  	       A  	           	       A  	       A  	       A  	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	           	           	       A  	       A  	           	       A  	           	       A  	           	       A  	           	       C  	       C  	       C  	       C  	           	       C  	       C  	           	   �� C  	           	           	       C  	           	           	       C  	       C  	       C  	           	       A  	       A  	           	       A  	       A  	       A  	           	       A  	           	       A  	       A  	           	           	       A  	       A  	           	       A  	       A  	       A  	       A  	       A  	       A  	       A  	           	       A  	       �  	           	       �  	       �  	       �  	       �  	           	       �  	       �  	       �  	       �  	           	       �  	       �  	           	       �  	       �  	       �  	           	       �  	           	       �  	       �  	       �  	           	           	       �  	           	           	       �  	       A  	           	       A  	   �� A  	           	           	       A  	           	       A  	           	       A  	       A  	       A  	       A  	       A  	       A  	       A  	           	       A  	           	       A  	           	       A  	           	       �  	           	       �  	           	       A  	       A  	           	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	           	       A  	       A  	       A  	           	       A  	           	       A  	       A  	           	       A  	           	       A  	   �� C  	           	           	       C  	           	       C  	           	       C  	           	       C  	           	       C  	           	   �� C  	           	           	       D  	       C  	           	       C  	           	       C  	                                   	       C  	           	       C  	           	       C  	           	   � C  	           	           	       C  	           	       C  	           	       C  	       C  	           	       C  	           	       C  	                                   	       C  	           	       C  	           	       C  	           	   � C  	           	           	       C  	           	       C  	           	       C  	       C  	           	       C  	           	       C  	                                   	       C  	           	       C  	           	       C  	           	   � C  	           	           	       C  	           	       C  	           	       C  	       C  	           	       C  	           	       C  	           	       P�  	           	       C  	           	       C  	           	       C  	           	   � C  	           	           	       C  	           	       C  	           	       C  	       C  	       C  	       C  	           	       C  	           	       C  	           	           	       C  	       C  	       C  	           	       C  	       C  	       C  	       C  	           	       C  	           	       C  	           	           	       C  	       C  	       C  	           	       C  	       C  	   �� C  	           	           	       C         C  	       C  	           	       C  	           	           	       C  	       C  	           	       C  	           	           	       C  	   /� C  	           	           	       C  	       C  	                  C  	       C  	           	       �  	           	           	       �  	       �  	           	       �  	           	           	       �  	   B� �  	           	           	       C                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      	       C  	           	       C  	           	       C  	       C  	       C  	           	       C  	           	       C  	           	       C  	           	       C  	   � �k  	           	           	   -� �k  	           	           	       �k  	   � �k  	           	           	       �k  	       �k  	           	       �k  	       �k  	           	       �k  	           	   �� �k  	           	           	   �� �k  	           	           	   4� �k  	           	           	   5� �k  	           	           	   C� �k  	           	           	       �k  	           	       �k  	       �k  	           	       �k  	           	   �� �k  	           	           	   �� �k  	           	           	   4� �k  	           	           	   5� �k  	           	           	   C� �k  	           	           	       �k  	           	       �k  	       �   	           	       �   	           	           	       �   	       �   	           	           	       �   	           	       �   	           	           	       �   	           	           	       �   	       �   	           	       �   	       �   	           	       �   	       �   	           	       �   	           	       �   	           	       �   	           	       �   	       @  	           	       @  	           	       @  	           	       @  	           	       @  	           	       @  	       @  	       @  	       @  	       @  	       @  	       @  	       @  	                       	       @  	       @  	       @  	           	       @  	       @  	       @  	           	       @  	       @  	           	       @  	           	       @  	       @  	           	       @  	           	       @  	           	       @  	           	       @  	       }   	       }   	           	       }   	           	       }   	       }   	           	       }   	           	       }   	           	       }   	          	           	          	           	          	           	          	           	          	           	          	          	           	          	          	           	          	           	         	           	           	          	           	          	           	        	           	           	          	          	           	    �    	           	           	          	           	          	           	   �    	           	           	          	           	           	       �   	           	       �   	           	    � �   	           	           	       �   	           	       �   	           	   � �   	           	           	       �   	       �   	           	    � �   	           	           	       �   	           	       �   	           	   � �   	           	           	       �   	       }   	           	       }   	       }   	           	       }   	       }   	           	       }   	           	    � }   	           	           	       }   	           	       }   	           	   � }   	           	           	       }   	       }   	           	    � }   	           	           	       }   	           	       }   	           	   � }   	           	           	       }   	           	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	      �   	           	           	       �   	           	       �   	           	     �   	           	           	       �   	       �   	           	    � �   	           	           	       �   	           	       �   	           	   � �   	           	           	       �   	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	       ]  	           	       ]  	   �� ]  	           	           	       ]  	       ]  	           	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	       ]  	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	   �� ]  	           	           	       ]  	       ]  	           	       ]  	           	       ]                                                                                                              	       c  	           	       c  	           	       c  	           	       c  	           	       c  	       c  	       c  	           	       c  	   �� c  	           	           	       c  	       c  	           	       c  	       c  	           	       c  	           	       c  	           	       c  	       c  	           	       f  	           	       c  	           	       c  	           	       c  	       c  	       c  	       c  	       c  	           	       c  	           	       c  	           	       c  	           	       c  	   �� c  	           	           	       c  	       c  	           	       c  	           	       c  	       c  	           	       c  	           	       c  	           	       c  	           	       c  	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	           	       m  	           	       m  	           	       m  	           	       m  	           	           	       m  	           	       m  	           	       m  	           	       m  	       m  	           	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	       m  	           	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	         	           	         	         	           	           	         	           	         	           	   �   	           	           	         	           	         	         	           	           	         	           	       m  	       m  	       m  	           	       m  	       m  	       m  	           	       m  	       m           	           	         	           	         	         	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	           	       ]  	           	       ]  	           	       ]  	           	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	           	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	           	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ^  	           	       ^  	       ^  	           	           	       ^  	           	       ^  	           	       ^  	           	       ^  	           	       ^  	           	       �  	           	       �  	       �  	           	           	       �  	           	       �  	           	   v�   	           	           	         	           	         	         	           	           	         	           	       ]  	       ]  	       ]  	           	       ]  	       ]  	       ]  	           	       ]  	       ]           	           	         	           	         	         	       ]  	           	       ]  	           	   �� ]  	           	           	       ]  	           	   �� ]  	           	           	       ]  	           	         	           	         	           	         	       ]  	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	         	         	           	         	           	         	           	         	           	   ��   	           	           	       �  	           	       �  	       �  	           	       �  	           	       ]  	       ]           	         	       ]  	           	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	       ]  	       ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       �  	           	       �  	           	       �  	       �  	       ]  	       ]  	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	                                                                                   	       �  	       �  	       :  	           	       :  	       :  	       :  	           	   ?� :  	           	           	       ;  	       ;  	       ;  	       ;  	           	       J  	       :  	       :  	       :  	       :  	           	       :  	       :  	       :  	           	       :  	       :  	           	       :  	       :  	       :  	       :  	       :  	           	       :  	           	       :  	           	       :  	           	       :  	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	   �� :  	           	           	       :  	   � :  	           	           	       :  	           	       :  	           	       :  	       :  	           	       :  	           	       :  	           	       :  	       :  	           	       :  	           	       :  	           	   �� :  	           	           	       ;  	       J  	           	       J  	           	       J  	           	       J  	           	   Q� J  	           	           	   �� J  	           	           	       J  	           	   �� J  	           	           	       K  	           	       K  	           	       K  	           	       K  	           	   8� K  	           	           	   �� K  	           	           	       K  	           	   �� K  	           	           	       L  	           	       L  	           	       L  	           	       L  	           	   g� L  	           	           	   �� L  	           	           	       L  	           	   �� L  	           	           	       M  	       �D  	           	       �D  	           	       �D  	           	       �D  	           	       �D  	           	       �D  	           	       �D  	           	       ^�  	       ^�  	           	       ^�  	           	       ^�  	           	       ^�  	           	       ^�  	           	       ^�  	           	       �D  	           	   �� �D  	           	           	       �D  	           	   �� �D  	           	           	       �D  	       �D  	           	       �D  	           	       �D  	           	       �D  	           	       �D  	           	       �D  	           	       �D  	           	   �� �D  	           	           	       �D  	           	   �� �D  	           	           	       �D  	       :  	           	       :  	                  :  	           	       :  	           	       K  	           	       K  	           	   �� K  	           	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	           	       :  	       :  	       :  	           	       :  	       :  	       :  	       :  	           	       :  	           	       :  	       :  	           	       :  	       :  	   �� :  	           	           	       :  	       :  	       :  	           	       :  	       A  	           	       A  	           	       A  	           	   � A  	           	           	       A  	       K  	           	       K  	           	       K  	           	       K  	                                                                                                                                                                       	       K  	           	       K  	       K  	       �  	           	       �  	           	       �  	           	       �  	           	       D  	           	       D  	           	       D  	           	       D  	       D  	       D  	       D  	       �  	           	       �  	       �  	       �  	           	       �  	           	       �  	           	       �  	                                                                                                                       	       �  	           	       �  	       �  	       C  	           	       C  	           	       C  	           	           	       C  	       C  	       C  	       C  	       C  	           	       C  	       @  	           	       @  	           	       @  	           	       @  	           	           	       @  	           	       @  	           	           	       @  	       @  	       @  	           	       @  	       @  	       @  	           	       @  	           	       @  	           	       @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	       J  	           	       J  	           	       J  	           	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	           	       J  	       J  	       J  	           	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	           	       J  	       J  	       J  	           	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	           	       J  	       J  	       J  	           	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	           	       J  	       J  	       J  	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	   �� J  	           	           	       K  	           	       K  	           	       K  	           	       K  	           	       K  	           	       K  	           	       K  	           	       K  	           	       K  	           	   �� K  	           	           	       L  	       J  	           	       J  	           	       J  	           	           	       J  	       J  	           	       J         �'             	       �'  	       �'  	           	       �'  	           	   �� �'  	           	           	       �'  	           	   �� �'  	           	           	       �'  	           	       �'  	           	       �'  	           	       �'  	           	   5� �'  	           	           	       �'  	           	       �'  	           	       �'  	           	       �'  	           	       �'  	           	       �'  	           	       �'  	           	   5� �'  	           	           	       �'  	       �'  	           	       �'         �             	       �  	       �  	           	       �  	           	   �� �  	           	           	       �  	           	   �� �  	           	           	       �  	           	       �  	           	       �  	           	       �  	           	   5� �  	           	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	   5� �  	           	           	       �  	       �  	           	       �  	          	           	   ��    	           	           	          	           	          	          	           	          	           	   ��    	           	           	          	           	           	          	          	           	          	           	          	           	          	           	           	          	          	           	          	           	   >�    	           	           	          	           	           	          	          	           	          	           	   ɝ    	           	           	          	           	           	          	          	           	          	       ]   	       ]   	       ]   	       ]   	       ]   	       ]   	           	           	       ]   	           	       ]   	           	       ]   	           	           	       ]   	           	       ]   	           	           	       ]   	           	       ]   	           	       ~   	           	       ~   	           	       ~   	           	       ~   	           	   Q� ]   	           	           	       ~   	       ~   	   D� ~   	           	           	       ~   	           	   E� ~   	           	           	       ~   	           	       ~   	           	           	       ~   	           	       ~   	           	       ~   	           	           	       ~   	           	           	       ~   	           	       ~   	           	       ~   	           	           	       ~   	           	                                                           
  _� ~   
  _� ~   
  �� �  
  �� �  
  �� D  
  �� D  
  4� K  
  4� K  
  D� ;  
  D� ;                                                                                                                                                                     ~                         	       ~   	           	       ~   	           	           	       ~   	           	       ~   	           	           	       ~   	           	       ~   	           	       ~   	           	           	       ~   	           	           	       ~   	       ~   	       ~   	           	       ~   	           	           	       ~   	           	       ~   	           	           	       ~   	           	       ~   	           	           	       ~   	           	           	       ~   	           	           	   Q� ~   	           	                  �             	       �  	           	       �  	           	           	       �  	           	       �  	           	           	       �  	           	           	       �  	       �  	           	       �  	           	       �  	           	           	       �  	           	       �  	       �  	           	           	       �  	           	       �  	           	           	       �  	           	           	       �  	       �  	           	       �  	           	       �  	           	       �  	           	           	       �  	           	           	       �  	           	           	       �  	           	           	       �  	           	           	       �  	           	       �  	           	           	       �  	           	       �  	           	           	       �  	           	           	       �  	           	           	       �  	           	           	       �  	       �  	       �  	           	   Q� �  	           	                  D  	       D  	       D  	           	       D  	       D  	       D  	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	           	       D  	       D  	           	       D  	   Q� D  	           	                  K             	       K  	           	       K  	           	       K  	           	           	       K  	       K  	       K  	           	   Q� K  	           	                  ;             	       ;  	           	           	       ;  	           	       ;  	           	           	   Q� ;  	           	              � ]   	           	           	       ]   	           	           	   n� ]   	           	           	       ]   	           	       ]   	           	       ]   	           	   � ]   	           	           	       ]   	           	    �  ]   	           	           	       ]   	       ]   	       ]   	       ]   	       ]   	       ]   	       ]   	           	       ]   	           	           	       ]   	           	       ]   	           	       ]   	           	       ]   	           	       ]   	           	           	       ]   	           	       ]   	           	       ]   	           	           	       ]   	           	           	       ]   	           	       ]   	           	       D  	           	           	       D  	           	       D  	           	       D  	           	       D  	           	       D  	           	           	       D  	           	           	       D  	           	           	       D  	           	    �  D  	           	           	       D  	           	   �  D  	           	           	       D  	           	    �  D  	           	           	       D  	           	   �  D  	           	           	       D  	           	    �  D  	           	           	       D  	           	   �  D  	           	           	   �� ]   	           	           	       ]   	           	       ]   	           	       ]   	       D  	           	           	       D  	           	       D  	           	           	       D  	           	       D  	           	           	       D  	           	       D  	           	       D  	       D  	           	       D  	           	    �  D  	           	           	       D  	           	       D  	           	       D  	           	       D  	           	           	       D  	           	           	       D  	           	           	       D  	           	   �  D  	           	           	       D  	           	    �  D  	           	           	       D  	           	   �  D  	           	           	       D  	           	    �  D  	           	           	       D  	           	   �  D  	           	           	       D  	       ]   	           	       ]   	           	       ]   	       |   	           	       |   	           	       |   	           	       �   	           	       |   	       |   	           	       |   	           	       |   	           	       |   	       ]   	           	       ]   	           	    �  ]   	           	           	   �  ]   	           	           	       ]   	       ]   	           	       ]          ]             	       ]  	           	       ]  	           	       ]  	                                               	   O� ]  	           	           	       ]  	           	       ]  	           	       ]  	           	   � B^  	           	           	   �� ]  	           	           	       ]  	           	       ]  	           	       �  	           	       �  	           	       �  	           	       ]  	           	       ]  	           	       ]  	           	       B  	           	       B  	           	       B  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	   Z� �k  	           	           	       ]  	           	       ]  	           	       ]  	           	   �� �   	           	           	       ]  	           	       ]  	           	           	       ]  	           	       �  	       �  	           	       �  	                                   	   ,� ]  	           	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	   �� ]  	           	           	       |  	           	   �� |  	           	           	       �  	           	       �  	                  |  	           	   �� |  	           	           	       |  	           	   �� �  	           	           	       �  	           	   N� �  	           	           	   6� |  	           	           	       n  	       n  	       n  	       n  	           	       n  	           	   �� n  	           	           	       n  	           	   6� {  	           	           	       n  	           	       n  	           	       n  	           	   �� n  	           	           	       n  	           	   N� �`  	           	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       |  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	                                                                                                                                                                                   	       ]  	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	       ]  	           	       ]  	       ]  	           	       ]  	           	   �� ]  	           	           	       ]  	           	   6� ]  	           	           	       h  	           	       h  	           	       h  	           	   �� h  	           	           	       h  	           	       h  	           	   �� h  	           	           	       h  	           	   N� m  	           	                  ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	                                   	       ]  	           	   �� ]  	           	           	   �� ]  	           	                  m  	           	       m  	           	       m  	           	   �� m  	           	           	   �� m  	           	                  �k  	           	       �k  	           	   	� �k  	           	           	       �k  	           	       �k  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	       �k  	           	       �k  	           	   �� �k  	           	           	       ]  	           	       ]  	           	       ]  	           	       ]  	                                                                                                                                                                                                                                                                                                                                                                                   	       ]  	           	       ]  	                                                                                                                                                                                                                                   	       ]  	           	       ]  	           	       ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	       ]  	           	       ]  	           	       ]  	           	       ]  	                                                                                                                                                                                                                                                                                                                                                                                   	       ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �I  	           	       �I  	           	       �I  	           	   �� �I  	           	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       /J  	           	       /J  	           	       /J  	           	       /J  	       /J  	           	       /J  	           	       /J  	           	       /J  	           	       /J  	           	   �� /J  	           	           	       /J  	           	       /J  	           	       /J  	           	       /J  	           	   r� /J  	           	           	       �I  	           	       �I  	       �I  	           	       �I  	           	       �I  	           	       �I  	           	   �� �I  	           	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	   r� �I  	           	                                                                       	   ��   	           	           	   �� n  	           	           	       n  	           	       n  	           	       n  	           	       n  	           	       n  	           	       n  	       n  	           	       n  	           	       n  	           	   a� n  	           	           	       �  	           	       �  	           	       �  	           	       �  	       �  	           	       �  	           	       �  	           	       �  	           	       �  	              �� �  	           	           	   |� �  	           	           	   �� �  	           	           	   �� �  	           	           	   i� �  	           	           	       �  	       �     �� �I  	           	           	   |� �I  	           	           	       �I  	           	       �I  	           	   �� �I  	           	           	   l� �I  	           	           	   i� �I  	           	           	       �I  	           	       �I  	           	       @J  	           	       @J  	           	           	       @J  	           	       @J  	           	           	       @J  	           	       @J  	           	           	       @J  	           	       @J  	           	           	       @J  	           	       @J  	           	       @J  	           	       @J  	           	       @J  	           	       CJ  	           	           	       CJ  	           	           	       CJ  	           	       CJ  	           	       CJ  	           	       CJ  	           	           	       CJ  	           	       CJ  	           	           	       CJ  	           	           	       CJ  	           	       CJ  	           	           	       @J  	           	           	       @J  	       @J  	           	       @J  	           	           	       @J  	       @J  	           	       @J  	           	           	       @J  	           	       @J  	       @J  	           	       @J  	           	       @J  	           	   �� @J  	           	           	       AJ  	           	       AJ  	           	       DJ  	           	       DJ  	           	       �J  	           	       �J  	           	       �J  	           	       �J  	           	       �J  	           	       �J  	           	   3� �J  	           	           	   d� �J  	           	           	       �I  	           	       �I  	           	           	       �I  	           	       �I  	           	           	       �I  	           	       �I  	           	           	       �I  	           	       �I  	           	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	           	       �I  	           	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	           	       �I  	           	       �I  	           	           	       �I  	           	           	       �I  	           	       �I  	           	           	       �I  	           	           	       �I  	       �I  	           	       �I  	           	           	       �I  	       �I  	           	       �I  	           	           	       �I  	           	       �I  	       �I  	           	       �I  	           	       �I  	           	   �� �I  	           	           	       �I  	           	       �I  	           	       �I  	           	       �I  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	   3� J  	           	                  J  	       J                                                                                                                                                                                                                                                                                                                                                                       	           	         	           	         	           	         	           	         	           	         	           	         	           	         	           	         	           	   ��   	           	           	   ��   	           	           	   ��   	           	           	   ��   	           	           	   |�   	           	           	   ��   	           	           	   ��   	           	           	   ��   	           	           	       4  	       4     �� ]  	           	           	   N� ]  	           	           	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	           	       ]  	       ]  	           	       ]  	           	       ]  	       ]  	       ]  	       ]  	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       n  	           	       n  	           	       {  	           	       {  	           	       {  	           	       �  	           	   .� �  	           	           	       ]  	           	       ]  	           	   1� ]  	           	           	       h  	           	       h  	           	       h  	           	       h  	           	       m  	           	       m  	           	       �  	           	       h  	           	       h  	           	       h  	           	       h  	           	       h  	           	       h  	           	       h         �  	           	       m         ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       n  	           	       n  	           	       n  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       h  	           	       h  	           	       h  	           	       h  	           	   e� h  	           	           	       �  	                  h  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       {  	           	       {  	           	       {  	           	       {  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	   �� �  	           	           	       �  	           	       �  	           	       �  	                  ]  	       ]  	           	       ]  	       ]  	           	       ]  	   �� ]  	           	           	   � ]  	           	           	       ]  	           	   �� �  	           	           	       �  	           	   � �  	           	           	   B� ]  	           	           	       ]  	           	   � ]  	           	           	       ]  	           	         	           	         	           	         	           	         	           	       i`  	           	       i`  	           	           	       i`  	           	       i`  	           	   1� i`  	           	           	   � i`  	           	           	   �� �  	           	           	   6� �  	           	           	   � �  	           	           	         	           	         	           	           	         	           	         	           	       � 	           	       � 	           	   �� �  	           	           	   � �  	           	           	   �   	           	           	         	   �   	           	           	       h  	           	       h  	           	       �  	           	       �  	           	       �  	       �  	           	       �  	           	       �  	       �  	       �  	       �  	       �  	           	       �  	           	       �  	           	       h  	       h  	       h  	           	       h  	           	       h  	           	       h  	           	       n  	       n  	       h  	       h  	           	       h  	                  h         ]  	       ]  	           	       ]  	       ]  	           	       ]  	         	           	         	           	         	           	         	           	         	                                                                                                                                               	         	   o� i`  	           	           	       i`  	           	       i`  	           	       i`  	           	       i`  	       i`  	         	           	         	           	         	           	         	           	         	           	         	           	           	         	         	         	           	         	           	           	         	         	         	         	         	           	         	           	           	         	           	         	           	   ��   	           	           	         	           	         	         	           	         	           	   ��   	           	           	         	           	         	         	           	         	           	   �   	           	           	         	           	         	           	   5�   	           	           	       �  	       �  	           	   � �  	           	           	       �  	       �  	           	       �  	       �  	       �  	       �  	           	       �  	       �  	           	       �  	           	           	       �  	       �  	           	       �  	                                               	       �  	           	       �  	           	       �  	       �  	   � �  	           	           	       �  	           	   � �  	           	           	       �  	           	       �  	           	           	       �  	       �  	           	       �  	           	       �  	                       	       �  	       �  	           	       �  	           	           	       �  	           	       �  	           	           	       �  	           	       �  	       �  	       �  	       �  	           	       �  	       �  	           	       �  	           	           	       �  	           	           	       �  	       �  	           	       �  	           	       �.  	           	       �.  	       �.  	           	       �.  	           	       �.  	           	       �.  	           	       �.  	           	       �.  	           	       �.  	           	       �.  	           	       �.                                                                                                                                                  	       �  	       �  	   � �  	           	           	       �  	           	   � �  	           	           	       �  	           	       �  	           	                                                                                               
  1� ?h  
  1� ?h  
  <� 4	  
  <� 4	  
  R� Cq  
  R� Cq  
  ]� �  
  ]� �  
  q� �O  
  q� �O                          
  �� �  
  �� �  
  j� �'  
  j� �'  
  �� �  
  �� �  
  G� ��  
  G� ��                                                                                                                                                                                                                                                                     ?h             	       ?h  	           	           	       ?h  	           	   � ?h  	           	           	       ?h         4	             	       4	  	           	           	       4	  	           	   ,� 4	  	           	           	       4	         ��             	       ��  	           	           	       ��  	           	   ,� ��  	           	           	       ��         Cq             	       Cq  	           	           	       Cq  	           	   �� Cq  	           	           	       Cq         �             	       �  	           	           	   R� �  	           	           	       �                                                                                                                                             �O             	       �O  	           	           	       �O  	           	       �O  	           	       �O                                                                                                                                 �             	       �  	           	           	       �  	           	       �  	           	       �  	                                                                                                           	       �  	           	       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	   �� ]  	           	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	       m  	           	   T� m  	           	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	       m  	           	   �� m  	           	           	       m  	           	         	           	         	           	         	           	         	           	         	           	         	           	         	           	       Ԗ  	           	       Ԗ  	                                                                                               	       m  	           	   �� m  	           	           	       m  	           	       m  	           	       m  	           	       {  	           	   �� {  	           	           	       {  	           	       m  	           	       m  	       {  	           	       {  	           	       {  	           	       �  	       �  	           	       �  	           	       �  	           	       �  	           	       �  	       �  	           	       �  	           	       �  	       �  	           	       �  	           	       �  	           	       �  	           	           	   �� �  	           	           	       {  	           	       {  	           	       |  	           	   �� |  	           	           	       |  	           	       |  	           	       |  	           	       |  	           	   �� |  	           	                  ]  	           	       ]  	           	       ]  	       n  	           	       n  	           	       n  	           	       �7  	           	       �7  	           	       �7  	           	       �7  	           	       �7  	           	       �7  	           	   T� �7  	           	           	       �7  	           	       �7  	           	       �7  	           	       �7  	                                   	       n  	       n  	       |  	           	       |  	           	       |  	           	       |  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	   �� �  	           	           	       �  	           	       �  	           	           	       �  	           	       �  	           	       �  	       �  	       |  	       |  	       m  	           	       m  	           	       m  	       m  	           	       m  	           	       m  	           	       m  	           	       m  	       �  	           	       �  	           	       �  	       �  	       v  	       v  	       �   	           	       �   	           	       �   	       �   	           	       �   	           	       �   	           	   T� �   	           	           	       �   	           	       �   	           	       �   	           	       �   	           	       �   	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	           	       J  	       �   	       �   	   w� �   	           	           	       �D  	       �D  	   $� �D  	           	                                                                                                                                                                                                                                                                                                                                                                                               	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	       ]  	           	       ]  	       ]  	           	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	   T� ]  	           	           	       ]  	           	   �� ]  	           	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	   �� ]  	           	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	   �� ]  	           	           	       ]  	           	       ]  	           	       ]  	           	       ]  	           	   �� ]  	           	           	       ]  	           	       ]  	       ]  	       ]  	           	       ]  	       ]  	           	       ]  	       ]  	           	       ]  	       ]  	           	       ]  	           	       ]  	           	       ]  	           	   �� �+  	           	           	       ]  	           	       ]  	           	   �� p- 	           	           	       ]  	           	       ]  	           	   � �  	           	           	       ]  	           	       ]         �+  	           	           	       �+  	           	       �+  	           	       �+  	           	       �+  	           	       �+  	           	       �+  	           	       �+  	           	       �+  	           	       �+  	           	       �+  	           	       �+  	           	       �+  	           	   7� �+  	           	           	   �� �+  	           	           	       �+  	           	       �+  	           	           	       �+  	           	       �+  	           	       �+  	           	       �+         p- 	           	           	       p- 	           	       p- 	           	       p- 	           	       p- 	           	       p- 	           	       p- 	                                                                       	   o� p- 	           	           	       p- 	           	       �S  	           	       �S  	           	       �S  	           	       �S  	           	       �S  	           	       �S  	           	       �S  	           	       �S  	           	       �S  	           	       �S  	           	   7� �S  	           	           	   �� �S  	           	           	       �S  	           	       �S  	           	           	       p- 	       p-        �  	           	       �  	           	       �  	           	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	       �  	       �  	           	       �  	       �  	           	       i  	       i  	           	       G  	       G  	   �� �  	           	           	   �� i  	           	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	       �  	       �  	       �  	           	   �� �  	           	           	       �  	           	           	       �  	           	       �  	           	       �  	           	           	       �  	       �  	           	   �� �  	           	           	       �  	           	           	       �  	           	   T� �  	           	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       <  	           	       <  	           	           	       <  	           	       <  	           	           	       <  	           	       <  	           	           	       <  	           	       <  	           	           	   �� <  	           	           	       <  	           	           	   �� <  	           	           	       <  	           	       <  	           	           	       �  	       �         �  	           	       �  	           	       �  	           	       �  	           	   p� �  	           	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	   �� �  	           	           	       �  	           	   7� �  	           	           	   ^� �  	           	           	   �� �  	           	           	       �  	           	       �  	           	       �  	           	           	       �  	           	       �  	           	       �  	           	           	       �  	           	       �  	           	       �  	           	       �  	       �         i  	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	   p� i  	           	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	   �� i  	           	           	       i  	           	   7� i  	           	           	   ^� i  	           	           	   �� i  	           	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	       i  	           	           	   �� i  	           	           	       i  	           	       i  	           	       i  	           	       i  	       i  	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	       �  	           	       �  	           	       �  	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	       �  	           	       �  	           	       �  	       �  	           	       �  	           	       �  	           	       �  	           	       �  	       �  	       �  	           	       �  	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	       �  	           	   3� �  	           	           	       �  	       <  	           	       <  	           	       <  	           	       <  	       <  	           	       <  	           	       <  	           	       �  	           	       <  	       h  	           	       h  	       h  	           	       h  	           	       h  	           	       h  	       h  	           	       �  	           	       �  	           	       �  	           	          	           	          	           	       w  	           	       w  	           	   � D�  	           	           	       w  	           	       w  	           	       w  	           	       w  	           	       w  	           	       w  	           	       w  	           	   	� w  	           	           	          	           	          	           	          	           	          	           	          	           	          	           	          	           	   	�    	           	           	       h  	           	       h  	       h  	           	       h  	           	       h  	           	       h  	       h  	           	       h  	           	       h  	           	       h  	           	       h  	           	       �  	           	       �  	           	   � �  	           	           	       �+  	           	       �+  	           	       �+  	           	       3  	           	       3  	           	       3  	           	       3  	           	   	� 3  	           	           	       h  	           	       h  	           	       h                    h                    h                    h                    h                �� h                               h         m         m         B^                    B^                    B^                    B^                    B^                    B^                 � B^                               B^                `� B^                           �� X^                           0� X^                           �� h^                               k^                    k^                �� k^                           �� k^                           �� k^                           C� �^                               �^                C� �^                               �^                    �^                C� �^                               �^                    �^                    �^                    �^                    �^                    �^                B� �^                           �� �^                           �� �^                               �^                .� �^                           �� �^                           �� �^                           �� �^                           �� �^                           �� �^                           �� �^                               �^                    �^         �                     �                     �                 �� �                             � �#                               �#                `� �#                           x� �#                           �� �#                           � �#                               �#                �� �#                               Р                    Р                    Р                    ��                    ��                �� ��                               Р                    Р         Р         Р                �� Р                               Р                    Р                    Р                    Р                5� Р                               ڠ         ڠ         ڠ         ڠ                0� 4�                           j� H�                           �� v�                               �                g� �                           �� �                           0� �                           �� )�                               ,�                    ,�                �� ,�                           �� ,�                           �� ,�                           �� F�                               Ģ                g� Ģ                           �� ٢                           x� ٢                           �� ٢                           �� �                               �                     �                     �                     �                     �                     �                                                                                                                                                                                                                                          � �                                �                     �                     �                 `� �                            �� �                            �� �                                �                     �                 4� �                                �                     �                     �                     �                 �� �                            �� �                            �� �                            �� �                            �� �                                :                    :                    :                    :                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    :                    :                    :                    :                    :                    :                    c                    c                    c                    c                    c                    c                    c                    c         c                    c                                                                                                                                                                                                                                                        :                    :                    :                    :                    :                    :                    �                    �                }� �                           ?� �                               :                    :                    :                    :                �� :                           ?� u                               c                    c         c         c         c         c                    c         c                �� c                               c                    c         c         c                    c                    c                    c                    c                    c                    c                5� c                               g                @� g                               �                    �         �                    �                    �                    �                    �                    �                    �                    �                    �                    �                    �                    �                    �                    �                    �                    �                    �                |� �                           �� �                           5� �                               �                @� �                               �                    �                5� �                           ��                                %                    %                    %                    %                    %                    %                    %                �� %                           �� %                               %                    %                4� %                               %                `� %                           �� :                           0� :                           �� J                               M                    M                �� M                           �� M                           �� M                           �� g                           �� �                               �                    �                �� �                           �� �                               �                    �                    �                    �                �� �                           �� �                           C� �                               �                C� �                               �                                                          ��                             �� �                               �         :                    :                �� :                           _� J                           �� J                           �� L                           C� L                               L                    L                    L                    L                    L                    L                    L                               L                               L                    L                               L                               L                    L                               L                               L                               L                           �� L                            � L                               L                    L                C� L                               L                    L                    L                    L                    L         L                    L         L                    L         L                    L         L                    L         L                    L         L                3� L                                                                                                                                                                                                                                                                                                                                                                                                                                                                               L                    L                    L                                                                                                                5� L                           �� M                                                                                                                                                                                                                                                                                                                                                                                           e                    e                �� e                           �� u                           �� u                               u                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         L                    L                    L                    L                    L                                                                    L                               L                               L                    L         L         L         L                    L         L         L         L                    L                               L         L                    L                               L         L                    L         L         L         L                    L                               L         L                    L                               L                    L         L         L         L                    L                               L                               L                                                                              � �D                               �D                    �D         �D                    �D         �D                    �D         �D                    �D         �D                `� �D                               �D         �D                    �D         �D                    �D         �D                    �D         �D                �� �D                           �� �D                           x� �D                           �� �D                           � �D                               �D                    D�                    D�                    D�                    D�                    D�                    D�                    D�                    A�                    A�                    A�                    A�                    A�                    D�                    D�                    D�         D�         D�         D�                B� D�                               D�                    ��         ��         ��                    ��                                                                                                                    ��                �� ��                               D�         D�         D�                    D�                �� D�                               D�         D�         D�                    D�                    D�                C� D�                               D�                P� M�                           �� �D                           b� g                               �                    ��                    ��                    ��                    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ��                    ��                    ��                                            ��                    ��                    ��                    ��                    ��                    ��                    ��                    ��                �� ��                           4� ��                           0� ��                           �� ��                           �� ��                               �                    �                    �                    �                                                                                                        �         �#                    �#                C� �#                               �#                    �#                    �#                    �#                    �#                    �#                ,� �#                           �� �#                               �#                    �#                    �#                    �#                    �#                    �#                    �#                    �#                    �#                    �#                    �#                    �#                    �#                    �#                    �#                    �#                    �#                �� �#                           N� �#                           �� �#                           5� �#                           � �#                               D�         D�         �#         �#         g                    g                C� g                               g                    g                    g                    g                    g                    g                ,� g                           �� g                               g                    g                    g                    g                    g                    g                    g                    g                    g                    g                    g                                                                    g                    g                    g                    g                    g                    g                �� g                           N� g                           �� g                           5� g                           b� h                               ��         ��         �         �         �                     �                 C� �                                �                     �                     �                     �                     �                     �                 ,� �                            �� �                                �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                                                                     �                     �                     �                     �                     �                     �                 �� �                            5� �                            �� �                                :     B� �                           �� �                           �� �                               �                .� �                           �� �                           �� �                           �� �                           �� �                           �� �                           �� �                           �� �                               �          �          �          �          �                     �                     �                     �          �                     �          �                     �          �                     �          �                     �          �                     �          �                     �          �          �          �          �          �          �         �         �         �         �         �                    �         �                    �         �                    �         �                    �         �                    �         �                    �         �                    �         �         �         �         �         �      �� �                            k� �                                �     0� �                               �          �          �                     �                     �          �          �                     �                     �                     �          �          �          �          �                     �          �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                     �                 |� �                            �� �                                �          �                     �                     �#                    �#         �#                    �#                �� �                            �� �                            �� �                            �� �                                �          :                    :                    :                    :                    :                    :                                                                                                                                                                                                                                                        :                    :                               :                               :                    :                               :         :                    :                               :         :                    :                    :                    :                               :                               :         :         :                    :         :         :                    :         �D                    �D                    �D                    �D                    �D                    �D                                                                                                        �D         �D         �D         �D         �D                    �D                               �D         �D                    �D                               �D                    �D                               �D                    �D                               �D                    �D                               �D                               �D                    �D                               �D                               �D                    �D                    �D                    �D                    �D                    �D                                                                                                        �D         �D         �D         �D         �D                    �D                               �D         �D                    �D                               �D                    �D                               �D                    �D                               �D                    �D                               �D                               �D                    �D                               �D                               �D         �#                    �#                               �#                               �#                    �#                               �#                    �#                               �#                    �#                               �#                               �#                    �#                               �#                    �#                               �#         �                    �                               �                               �                               �                               �                               �                               �         �                 o� �                                �                                �          �                     �                     �                     �                     �                     �                     �                     �                     �                     �          �                    �                    �                �� �                               �         �                                                                                                                                                                                                   ��                                                  �         �         �                    �         �                    �                �� �                               �         �         �         �                                                                                                                                                                                                                                                                                 ?h         ?h                    ?h                                                                                ?h                    ?h                                            ?h                �� ?h                               ?h         4	         4	                    4	                                                                                4	                    4	                    P�                    4	                �� 4	                               4	         D�                    D�                    D�         D�                    D�                    D�                �� D�                               D�         D�         �                �� �                               �         �                                                                                                                                                                                                                                                                                 i`                    i`                                    ��                                                  i`         i`         ]                    ]                    ]                    �         ]                    ]                    ]                                                        ]                    ]         ]         ]                    ]                    ]         ]                    ]                    ]                    ]         ]         ]         ]         ]                    ]         ]                    ]                    ]                    ]                    ]                    ]                �� ]                               ]                    ]                    `                    `                    `                    `                    `                �� �i                           �� �i                           �� c                           �� c                           �� ]                           �� ]                           .� `                           �� `                           � Ci                           �� ]                               ]                    ]                    ]         ]                    ]                    ]                    ]         ]                    ]                    ]                    ]                    ]                    ]                    ]         ]                    ]                    ]                    _                    ]                    ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ]                    ]                    ]                               ]         ]                    ]         ]                    ]                               ]                    ]         ]                    ]         ]                    ]                    ]                    ]                    ]                    ]                    ]         ]                    ]                    q                d� q                               q         q         q         q         q                    q                d� q                               q                �� q                               ]                    ]                    ]                    ]         ]                    ]                    ]                    ]                    ]                |� ]                               ]                :� ]                               ]                    �         ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]         ]                    ]                    ]                    ]                    ]         ]         ]         ]                    ]                    ]                                                                                                                    ]                    ]                    ]                    ]                    ]                    ]                    ]                0� ]                               `                    ]                    `                    `                    `                    `                    `                    `         `                    `                    `         ]                    ]                    ]                    �                    �                    �                    ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     c                    c                    c                    c                                            c         c     �� c                               c                �� c                               c                    c                          �� c    �� c    i� �    i� �    �� c    �� c    �� �    �� �    v� w    v� w    �� �:    �� �:    *� (    *� (    o� h    o� h                                 �i                    �i                    �i                    �i                �� Wn                               Wn                � Wn                           �� �                               �                � �                               �i                    �i         �i                                                                                                                                �i                    �i                    �i                    �g                    �g                    �g                    �g                    �g                    �g                    �g                y� �i                               �i         c                    c                    c                    c                    c                    c                    c                    c                    f                    f                �� f                               f                d� f                               f         f                    f                    f                d� f                               f         f                    h                    h                    h                    c                    c         c         c                p� c                               c                    c                    c                    c                    c                    c                �� h                               h                    c                    c                �� c                               c                � g                           ]� g                           �� }                               }                � c                           y� c                           � c                               c         c                �� c                               �                    �                    �                �� �                               �                    �                    �         �                p� �                           � �                               �                �                            ��                            � �                           � �                           �� �                               c                    c                    c                �� f                               c                    c                �� ��                               ��                                                        c                    c                    c         c                p� c                           �� c                               c                    c                3� c                               c                    c                    c                    f                3� f                               f                � c                           �� c                           � f                           y� c                           � c                           �� c                               �                    �                    �                    �                    �                    �                    �                    �                    �                    �                    �                    �                T� �                               �                    �                    �                    �                    �         �                    �                    �                    �                    �                    �                    �                    �                    �                    �                    �                    �         �                    �                    �                    �                    �                    �                ;� �                           �                                                                                        ;�                                �                    �                    �                    .                    .                � .                               �                    �                    �         �                p� �                               �                    �                    �                    �                    �                    �                ��                                                    �                    �                �� �                               �                �                            m�                            �� G                               G                � �                           y� �                           � �                           �� �                               w                    w                    w                    w                    w                    w                S� z                               w                    w                    w         w                p� w                           � w                               w                �� �                               �                � �                           �� �                           � w                           � w                           �� w                               �:                    �:                    �:                    �:                    �:                    �:                    �:                    �:                    �:                    �:                �� �:                               �:                    �8                    �8                �� �8                               �:                    �:                    �:                �� �:                           �� �:                               �:                    �:                    �:                    �:         �:                p� �:                           �� �:                               �:                �� �:                               �:                � �:                               �                    �                    �                y� �                               �                    �                �� �                           � �                               �                    �     y� �                               �         �                    �                    �                $� �                           � �:                           $� �:                           ��  �                                �                �  �                           $�  �                           � �:                           � �:                           �� �:                               (                    (                �� e5                               (                ]� (                               (                    (                ]� (                               (                    (                ]� (                               (                    (                ]� (                               (                    (                    (                    (                    (                    (                    (         b5                    b5                    b5         (                p� (                           �� (                           |� (                               (                6� b5                               b5         (         h                    h                    h                �� h                               h                    h                    h         h                p� h                           � h                               h                    �h                    �h                � �h                           �� �h                           � h                           � h                           �� h                               �m                    �m                    �m                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     �:                    �:                    �:                    �:                    �:                    �:                    �:         �:                    �:                T� �:                               �:                �� �:                               �:                    �:                    �:                    �:                �� �:                               �:                    �:         ��         ��                                                                                                                                                                                                                                                                                                             d�                                                             D                    D                    D                R� D                               �                d� �                               �         �                    �                    �                             z                    z                    z                    z                    z                    z                �� z                               z                    z                    z                    z         z                    z         z                    z         z                �� z                               z                    z                    z                    z         z                    z                    z                    ��                    z         z                    z                    z                    z                    z         f                    f                    f                    f                    f                    f                    f         �                d� �                               �     �� �                               �                    �         f                d� f                               f         f     �� f                               f                    f         m         �#         h         �         f         z         ��         ��         }                    }         }         }                    }                �� }                               }                    }         �                    �                    �                �� �                               �                    �         �#                    �#                    �#         h                    h                    h                    h         h                    h         h         h                    h         h                    h                �� h                               h                    h         s                    s                    s                �� s                               s                    s         z                �� z                               z         c                    c                    c                    c                    c                    c                    c         f                    f                    f                    f                    f                    f         Ci                    Ci                    Ci                    Ci                               Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci                    Ci         Ci                    Ci                �� Ci                           � Ci                               Ci                    Ci                    Ci                    Ci         Xi                    Xi                    Xi                    Xi                    Xi                    Xi         [i                    [i                    [i         [i         [i                    [i                �� [i                           � [i                               [i                    [i                    [i                    [i         �i                    �i                    �i                    �i                    �i         �i                    �i                    �i                    �i                    �i                    �i                    �i                    3	                d� 3	                               3	                    3	                         ��                            ��                                3	                    3	                    3	                    3	                    3	         3	                    3	                    3	                �� 3	                                                                               3	                    �i         �i         �i                    �i                    �i         �i         �i         �i                    �i                    �i                    �i                    �i                    �i                    �i                    �i                    �i                    �i                    �i                y� �i                               �i                     |         Bq         kx         �                  �O                     �         c         c                    c                    c                    c                    c                    c                    c                    c                    h         h                    h                    c                    c                    f         f                    f         f                    f                    f         f         f         f         f         f                    f                    f                    c         c                    c                    c                    c         c     3� c                               c                4� c                               c                    c                          ;� e5    ;� e5    K� e    K� e    q� c    q� c    �� �:    �� �:         e5                    e5                    e5                    e5                    e5         -�                    -�                    -�                    -�         e                    e                    h                    h                    h                    �                    h                    h                    h                    h                    h                    e                    e                    e                    e                    e         n                    n                    n                    n         c                    c                    f                    f                    f                    i                    f                    f                    f                    f                    f                    f                    f                    f                �� f                               c                    c                    h                    h                    h                    h                    c                    c                    c                    c                    c         l                    l                    l                    l                    l                    l                    l         q                    q                    q                    q         �:                    �:                    �:                    �:                    �:                    �:                    �:                    �:                    �:                    �:                    �:                    �:                    �:                    �:                    �:         �:                    �:                    �:                    �:                    �:                    �:         c                    c     �� c                           � c                               c                    c                    c         c                |� c                               c                6�                            :� c                               c                    g                    g                    s                    �         �         s         s                    s                � s                               ^                    ^                    ^                    ^                    g         c         c                    c     �� �                           |� �                               �                6� j\                               j\         j\     � �                               �                                                                                                    �                                                                                                                                                                                                                                                                                                                                                                                                                              ��                                                                                                                                                                                                                                                                                                             c                    c                    c                    c                    c                    c                    c                    c                    c                    c         c                    �                    �                    �g                    �                �� �                               c                    c                    c                    c         c                |� c                               c                T� c                               c                    c                    c                    c                    c                    c                    c         c                    c                    c                    c                3� c                               c                    z                    z                    �                3� �                               �                    z                    z         z         c                    c                    c                    �         �                    �                    c                    c                    c         c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             c                    c                    c                    c         ]                    ]                    ]                    ]                T� ]                               ]                �� ]                               ]                    ]                    ]                    f                �� f                               f                    ]                    ]                    ]                    ]                    ]                    h                �� h                               h                    h                    h                    m                �� m                               m                    ]         ]                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ]                    ]                    ]                    ]         z                    z                    z                    z                    �                    �                    �                    �                    �                    �                    �                    �                G� a                               �                    �                    �                    �                    �                C� �                               �a                    �a                    �a                    �a                    �a                C� �a                               z                    z                    z                    z                    z                    ^                    ^                    ^                    ^                G� :                               ^                    ^                    ^                    ^                    ^                    ^                    ^                C� ^                               �                    �                    �                    �                    �                    �                    �                �� ^                               ^         z         z                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]                    �                    �                d� �                           K� �                           �� �                               ]                    ]         ]                    ]                    ]                    ]                    ]                    ]                    ]                    ]         ]                    ]                    ]                    ]     �� �                               �                    �                    �                    �                    �                    �                    �                    �                    �                p� �                           @� �                           � �                               �                �� �                               �                    �                    �                    �                    �                    �                    �                g� �                               �                    �                                                    Q� �                               �                    �                �� D                               �                    �                    �                    �                    �                    �         �                    �                5� �                           �� �                               �                    �                �� �                           � �                               �                �� �                               �                    �                    �                    �                                                                                                                                                                                                                                                                                                                    �                               �         �                    �                    �                    �                    �                    �                    �                    �         �                               �                               �         �                    �                               �                    e�                    e�                               e�                    e�                           � e�                               �                    �                )� �                               {                    {                5� {                               �                    �                    �                    �                    �                    �                    �                    �                s� �                           �� �                               �         �                    �                    �                    �                    �                    �                    �                    �                    �         �         �         �                    �                    �                    �                    �         �         �                    �         �                    �         �                    �                    �         �         �         �         �         �                    �                    �                    �         �                    �                    �                    �                    �                    �                    �                    �         ]                               ]                    ]         <                    <                    <                    <                �� <                               <                    <                    J                    J                    J                    �                    �                    �                    �                                                                                J                    J                    J                    J                                                        J                    J                    J                    J                T� J                               J                    J                    J                    J                    J         J                    J                    J                                                                    J                    J                    J         J                    J                    J                    J                    J         J         J                    J         J                    J                    J                    J                    J                    J                3� J                           �� K                               <                    <                    <                    <                    <                    <                    >                    >                    >                �� <                               �                    �                �� �                           � �                               �                :� �                               �                |� �                               �                �� �                               �                    Ai                    Ai                    Ai                               �                    �                    �                    �                    �                    �                    �                    �                �� �                                                                                           !i                    !i                    !i                    !i                                                                                                                                                                    �                    �                    i                    i                    i                    i                    i         i                    i                    i                    i                    i                    i                    i                    i                    i         i         i                    i                    i                    i                    i                �� i                               �                    �                    �                    �                                                                            �� �                           �� <                               <     t� ]                                ]                     ]                 `� ]                                ]                     ]                     C^                    C^                    C^                    I^                    I^                    I^                    I^                               C^                    C^                    C^                    C^                               C^                    C^                               C^                    C^                           �� C^                           �� ]                                ]                     ]                 �� ]                                ]                     ]                 n� ]                                ]                     ]                 	� ]                                ]                     ]                 � ]                            �� ]                                ]          ]                     ]                 ^�                                 ]                     ]                 H� ]                                �                     �                     �                     �          �                     �                     I     �� I                           �� I                           �� �                           ^� �                           k� �                                �                     �                     �          �                 �� �                                �                     �                     �                     �                     �                                �                     �                                �                     �                     �                     �                            �� �                            H� �                            �� �                           H� �                               ]                     ]          ]                               ]                     ]                 � b                                b                            E� ]                                ]                     ]                                                                                                                                                                                  ]                     ]                                      ��                                             ]                     ]                 �� ]                                �                     �                     �                     �          �                     �                     �     �� �                           � �                           �� �                           �� �                           k� �                                �                     �                     �          �                     �                     �                 k� k                           �� k                           �� �                                �                     �                     �                     �                     �                                �                     �                                �                     �                                �                     �                     �                     �                            �� �                            �� �                                �                    �                    k     �� �                           �� �                               ]                     ]                     ^         ]                     ]                     ]                     n         ]                     ]                 � b                                b                            E� ]                                ]                     ]                                                                                                                                                                                  ]                     ]                 T�                                 ]                     ]                     ]          i                     i                     i                     i          i                     i                     �     �� �                           � �                           �� �                           T� �                           k� i                                i                     i                     i          i                 �� i                                i                     i                     i                     i                     i                                i                     i                                i                     i                     i                     i                                i          M                    M                               M                    M                    M                    M         ]                     ]                     ^                    ^                    �                    �                    �                    �                    �                    �                    ]                     ]                     ]          ^                    ^                    ^                    ^         ^     @ ^                               ^                @ ^                               ^                    ^                    ^                    ^                    ^                    ^                    ^                    ^                    ^                �� ^                               _                    _                �� _                               ^                    ^                    ^                    ^         ^                    ^                    ^     �� ^                           �� ^                               n                    n                    n                    n                    n                    n                � n                           k� ^                               ^                    ^                    ^         ^                �� ^                               ^                    ^                    ^                    ^                    ^                               ^                    ^                               ^                    ^                    ^                    ^                           �� ^                           �� ^                           �� �                           �� �                               ^                    ^                    ^                    б         ^                    ^                � ^                               ^                           E� ^                               ^                    ^         n                    n                    n                    n                               n                    n                    n                    n         ]                     ]                 ��                                 ]                     ]                 k� ]                                i                     i                     i                     i          i                     i                     �     �� �                           -� �                           �� �                           �� �                           k� i                                i                     i                     i          i                     �                    �                    �                    �                    �                               �                    �                           �� �                           k� �                           �� i                            k� i                                ]                     ]                     ]                     ]          �                    �                � �                               �                           E� �                               �                    �         �                    �                               �                    �                    �                    �         �                k� �                               �                    �                k� �                               �                    �                k� �                               �                    �                    �                                �         �     �� �                               �                �� �                               �                    �                    �                    �                          �� �    �� �    �� �    �� �                            � I    � I    � �    � �         �         �                    �         �         �                    �                    �                    �                    �                    �         �         �         �         �         �                    �     �� �                               �                    �         �                    �                    �                    �                    �                    �                    �         �                    �         �                    �                    J                    �         �         �                    �                    �                                             I                    I         �                    �         A                    A                    A                    A                    �                     A                    A         A                �� A                               A                    A                    A                    A                    A                    A                    A                    �          �                     A         A      @ A                               A                @ A                               A                    A                    A                    A                    A                    A                    A                    A                    A                    A         A                    A         A                    A                    A                    A                    A                    A                    A                    A                    A                    A         A                    A         A                    A                    A                    A                    A                    A                    A         A                    A                    A                    A                    A                    A                    A         A                � A                               A         i                     i                 k� i                                i          i                     i          i      �� i                                i                 �� i                                i                     i                     i                     i          i                     i                     i                     Y                    i          i          i          i          i          i                     i          i                     i                     i          i                     i          b                     b          b          b                     b          b                     b          b          b          b          b                     b          �                     �                     �                 �� �                                �                 �� �                                �                 �� �                                �                 �� �                                �                     �          i                     i                     i          i                     i          i                 �� i                                i                 �� i                                i                 �� i                                i                     i          �                    �                    �                    �                    �                    �                    �                    �                    �                                                                                             b                     b                 �� b                                b                     b                     b                     �          �                     �                     �                                                                                 b          b                     b                     b                     �                     b                     b                     b                 �� b                                b                     b                     b                     b                     b          ]                     ]                     ]                     �                     �                     �                     �                     �                     �                     �          �                 �� �                                �                 �� �                                �                 �� �                                �                     ]          ]          i                     i                     i                     I                    i          ]                     ]                  �  ]                            �  ]                                ]          ]       @ ]                            @ ]                                ]          ]                  @ ]                                ]                 @ ]                                ]                  @ ]                                ]                 @ ]                                ]          ]                  @ ]                                ]                 @ ]                                ]                  �  ]                                ]                 �  ]                                ]          i         i         �          �          �          �          �         �         �          �          ;         ;         )         )         �          �          i          i          �         �         A         A         f         f         �         �         I         I         I         I         I         I         I         I         J         J         J                     i          i          i                                                                                                                                                                                                                      �         �         �         �         �         �         �         �         �         �         �                     �         �         �                                                                                                                                    {         {         {                     ^         ^         ^         ^                                             ^                                                         �         �         �                     �          �          �          �          �          �          �          �         �          b          �                      �         �         �                                                                                                                                                                                                                                                                                                                                                                                                                     >         >         >         >         >         >         >         >         ?         ?         ?                     >         >         >                     �          �          �          �          �          �          �          �          �          �          �                      �          �          �                                                                                                                                                                                                                      G         G         G         G         G         G         G         G         H         H         H                     �         �         �                     c         c         i         i         ]         ]                                 h         h         �#         �#         z         z                                 (         (         ��         ��         z         z                                                                                                                                                         �         �         �         �                                 K         K                                                                                                                                                                                                                                                                                 B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         B         @         @         @         @         �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          �          A         A         A         A         m         m         m         m         e�         e�         e�         e�         �         �         �         �         �A         �A         �A         �A                                                                                                         B         :         C         C         C         C         o         o         o         o         g�         g�         g�         g�         �         �         �         �         �A         �A         �A         �A                                                                                                                                                                                        �                              �                                                                                                                                                                ��       ��       ��       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         